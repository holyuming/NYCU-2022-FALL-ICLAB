`include "../00_TESTBED/pseudo_DRAM.sv"
`include "Usertype_FD.sv"
`define CYCLE_TIME 3.2
`define PAT_NUM 200*10000
`define THRESHOLD 100

program automatic PATTERN(input clk, INF.PATTERN inf);
import usertype::*;

class random_data;
    rand Action action;
    rand Delivery_man_id deliver_id;
    rand Ctm_Info cust_info;
    rand Restaurant_id rest_id;
    rand food_ID_servings food;

	constraint limit {
        action dist{Take:=3, Deliver:=2, Order:=2, Cancel:=5, last_data.action:=5};
		deliver_id dist{[0:255]:=1, last_data.deliver_id:=255};
        cust_info.ctm_status inside{2'b01, 2'b11};
        cust_info.res_ID inside{[0:255]};
        cust_info.food_ID inside{[1:3]};
        cust_info.ser_food inside{[1:10]};
        rest_id dist{[0:255]:=1, last_data.rest_id:=255};
        food.d_food_ID inside{[1:3]};
        if (action == Cancel)
            food.d_ser_food == 0;
        else
            food.d_ser_food inside{[1:15]};
	}
endclass

//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
fYP110p9zIKGg9jvB1QSdBIGlIiFvYNUW9sKnbr/h80nUY47P8i7uwUCixvml+Eq
c9d98uN2eXYuRcTq3OYSSJ/QKjJ7wbHRw8ZZZqRIN5or6Kt6fUM7xEff9S92Hf4r
lQy284R+Bpi/lWE0WvNO/K6zdHiMrOQZMWTpRgTln9qRs6u2v7l8seH0Q95dIjKg
na6B6y/HZs7BEcVaTpaLJoT7S2hKLrt6lIRK77MBKZ5zrAlmPy8o1rtjJIOhFkvx
wLOzDnbFtjRvQQNGv2DmFEirvqmdlNLHaQnVzEaBKDW5S91v0OV+XnbHFPjpk58E
oY6hm7Sobu5ErpV1JqvShA==
//pragma protect end_key_block
//pragma protect digest_block
L+W8F5amH8e0Pdh5myRi+Wir54k=
//pragma protect end_digest_block
//pragma protect data_block
SmtfHdtkeqF7zz7fv1j0g3/LwW8/7UC/O7Cu8Jk+xK6XsluHtqIiXoDTJ0vquwDU
s3tAQ5AhArPWs1BSY2ZG2Q61EGjQaj2fluYVt1EBfdhwMy4/1ToQRqRkddt+4uu0
1rej5FxpMUYfq8giib1RLP6k14dOonitwjXECH6BGdFBhA4Y3EvL3n/nAm3vvLKp
46UNn2XwLD9yx0L3hCZljs/kijSRCDqHzBHLrBjP1UlvesV+GNxn1iW7ClsoWFyC
+THfnICiJFQ4BWmuhxhW39kVRElrWzuC4WEnzkwAmo6oMZPp9dwvJJlAKySV2ZiL
BzqaZMcvn/bE++jmeXHEgZTzgFnVFop+CR3KnRjZ23IL/FhoCTLdMOt5ULb/rctv
SHhMptX47xJ8wsbKOVQURijF0JB42B3HQv3CyxeigmFNDMaMjFqaa3NjRLXUy/Lz
ujJJE73HF60Vqz+2+/Vv8FPq4fxWTkHlAJNfCWA22PqK4BYOm/tM9R9CLORFHLoL
PL6ELNB5DjTwYZfNeNrqXXKMf40Aoo33c8J5rbdUEAXipPrHx8swY3N9rlv5uMJE
aMDaijalOB29YSFsRThQh0sA5kVtTTiXqvbAjtT9YWWX0l5KhHXCiaotOJPjAOY+
hbbcNCxGcmxSWT48M87/4LuxU3bFAfVJ6GEBLaEU2nPjKocKySEk9G7pAW0/CM6p
5+q2i8tkwJj3MKI+ASgopCrQ6AeOzeA9+4qv2zn5IY++yYdQenKNXLGAh+n209Ue
AE/fS8pGYEEXp6eK05AmIVZRMXSekEjMOgjYC++THX7qxGxDaWheew/m5Ks0PROB
MEpv/3B/A/5WNfHBOsx83EDqfEabl7Lh9jq99MkEezXY0aJX8u2dvtH3fwhKLF/0
22byceKW5aB6dLqrmH4tbbst/BUC4hwVKN+mj8c5pBPI442oy2WqMokbBOORqZZb
KUf+I1BJd5GX/ELa20/BL8vUpfhqz9Yb3zgjSGusxpM4rWQfb9CoAb9AZQDr8Q11
ZueBdeoQCM99fvZjjnzlaPLLUV0OTCmsbheeroNMCBUxZmVx9mLuUn00W6y90akC
jaSvQ3mtMaeDbXa0gM6k+s52fghLC0nOYGP7hc72qZuE2a+PoUKi4pA/3aCl6RTS
dHMjm7EQYmUSjQKxn0BqKERLefdx7HR4noAvQHcZYVTmLAhqrrfXHUgm2oxazsBp
edji6ckNwz8W3n2FJtvQNmvjnN3DBZgFA1//Xwyf+3VjAnHSxW8Cv9I9tqxayTGB
bmSt5Sbg08rY2uN6kT0NAt7Gr3IXtk7iRwQORfR1OyGtLlbtVPxGsqGmTG6VVMkt
Ve5p9d/M83UUtplP797q/7fb8FuI+AMmmqTTVFy6ubJulOSG2ToPAYViKGVQmpaI
ACqTWWMBsFkeaEnNAmTWWBVhbPK9x3VLZ0fr4Q/COLmOpUpcNmmUtsqN/MSvIVIY
ZUANA8Ow4XzRD8UGWtXieVXK3AukpqJ+bMysemepvrEGL4MSn+kT9XtUXIV3wKQd
nks7Hzh9oFlrbW/RMs6KGobOP7QdBuWuQZnTLqVMv9rhunRpqFQqULrXoxezmQLo
i6jCsVVDgp63zaalSn1p26bNLgyCB7Uifi0HNB0WNADLFsLm3BNgLds2DBOXLq8s
Ctq5pQdSdHNnS+rohWP8S4gbNr6SWO4q/UDt4TO0OxVDe0/iUoYG41nX7Q4HhfOA
62Mk5IrsiPuFwqlt1dGzPGM2FuDALPg4O/OateNdNInPRkMcJMalG/mnhzV8Vu01
9SE8sm2bG3DmL6zRfCSPNA3j2JzhfAFP5mUluPM1+ShP7fUAxNOfQzV7OBPlIRJA
H5C2WlYypgYEz/jVG/A+ep7AawNBACNZ+7yl8cWLo/WexqdBaLMp/YFFqlm3bf0B
ZBS2Ufh+zf5EgFHyLWZlx02zKPYqI9u6L4a5CZ4SWE16FNQI7eVvW/jH2ecsz1Sw
Dm4ZkW2mYFEB3FbEMui/5fk++d/+h82pzuwCs7ZKM77ZTWOzTakNLP4STyLrDfQu
/BhMTKeoMOTmxtecDkuxvTTpS+Fse+Gyd6vRrTrj0wkQ1y3jMIjZpMq6DnsPBwp3
7BMYzzT/2j+UYn9eHjWOf/ierLYWxg01Vaff+sOm85flqotdzLrX/0KOUnbVr+RE
e90DZtQHeufupKrSqOph4oBMQB3oZXd23QyKFISnUrbNRHgqZUlpgVgAqpMOjwZY
rZ2vpyw07WDw+raLaJn/IsANtDmZxQHdBnhR6EQkM5OszAYeVQd2EqdTFEhu4tKc
ijLfvPALf1FzoY0Rb4lagia4g0zoWwtjeLhTyW9ARNoUiwLdxKUSLaePMZVx/a+8
EzrT2kv8MIm9x1+/ZwqtdEItHIHQc++H8/1LlcRJBEs+zlJaD5OGaWwlNvX92ny3
wC6vKSXYDcWlZzBRQPgWl57hv+HII+zzrEif5yNfkzZ1SpLAQjANbO00bURqBJ5o
Go3LRoXD63kS3r3LHPncRulG4iLccywkiXHzul8UQ5kKQoUU2t9NoUGSkrU3WzEs
TXY3hmGvvIQpTESm+obUBuFFkos3VI190MXq6yJR+ry+sx+mFJfsVx1+H0x9rza2
atqcOHvsWSNFqkHA3mxu5AjIsKhho4MFBES9A7BJN0UfabBLQiDR4KRC5LTq6t8C
GcAvZ/btFvb1h1rU0xr8xV8hmuQB/jcbNOddcD7GpMfIG0RkoPkBB94/g6QBEjfZ
fdsVwz7Ds0NOWvvqyLclbvP/VU1I33IsngtDUbNIib2JfvdJUKfnMWq7d7Zmk5zS
dzj6ygEStkGVcxzZHDCWka7Z7iCXxLpTRb6yLgPdD6AyLpj5Y2tMPY8Yi7vdx4rs
6xelmAoaqNRcHrpx+r3a95zvVDTRGLEQE8cx/UDzVcl4+mMXGtN+MapNlgFKramm
1syV8RuBbaD4x5RHMBrKrv5u3t0G0S83RpmOOX1rvJy19yG4UASV08IqnENbuetJ
Ch2koOZJTozhaxksUMXbAB5ONKxHlGS14HnUQ6XILOygEns7S5to3emJIEYkX7Wy
cyL4Dzzcr8HkvkT9IQ3ISUDKmDSZc40yIfMAuh+giBRUs6yNtI4q+oby36LsgfC6
pV+GoDPcwV66AnDV73k+I1wrO6lX9RkdUdPAUykFOa0iaLyYzb5NjWkxr5/SA6hE
9uZHTDaeETNIQncYiZVlomLTHuHgVJI//uas4eMMABFMIaYPvfm4gqnvsBzK6Lcm
p37URfDWvhC3JaUwqcx8CP/HJcCWdUbpC7upkdr5HxiHGxQYrPFgYtj12lbJKDM8
HujQXSShcKZCST2ETRw73HUqzBcCBrFmhrgZs3bVRVbopi6xlYiq+EvZaDWK1v6Z
gPPJWwT+FT2a8B70B8Q/VsHWBzAh4GY1oh/pENqKUFxP1vK+1wN7asTvSGGfMJ5J
miGDyaV8vAmQnvMYDK2p03syxUPca2K8rYZXSzVxJpfDqh8IY26XGev+PGRKA/WU
Nxr3++G9hifaQsYb//uC7U8oAzJcAqxsOndQnW+jHloqbb2RjdWaoAjRRJ/nmxiI
89h3tXFnpYxFgJhoUd++N3d2s5LcpZA2hh4uOo52fergu+hRbuomsgL6F4bHQNyw
GZVKZYn4mguW8Nw320Yqv16lTTlh+ThaFc4JGGQXvHbzfjRz0v8cXQmgnWHxHtSR
FcYhCMGoDH9U5KhV1xSHqlq/MEjkY4DpM3XE5F4ZOJVOaUIUQeJC03ReOJkZM3i2
PvpjoGkU8UUONZ6m5g84dRDf+Stegt0xzhCUsPE5IdFgjtC51B+mUaq/pFrKgqgy
JZcAFsBTcTL74W/DSSMFV1m8sw5nqRnkvKzBc0ALzRhsb/KsOEiW9ZarhIyatvuE
+m/gLvWOwQ6aWiubApTrMPMOvO81gEPQHfYg12DALorfvRnK2kVOwpxy+UayRLhS
7IWw+lfQKsz6/F0hHyCQd3L4rkdXO7hHLCZNX+Cq77w26y7/WFzms3afHMeg0OP3
szlJ9Wojp41TPj0qtds8yxLZ7DKRsPWf6OPQStcuydpGHCztyDxShn+hJieSOnz+
GgJQ4tkcCRAroDnyOMZuZIqnnPDn44hr12FNJ2g9Dtmi9ZlJ77s8fnCRqaUdd0W5
mpCuhf9XjH1YU1NNVAOsOCXuQ+xmzm/zPOPUbgSzxvKd39CRPLeXOsi4IpdIZPRf
OLaSfAjYSG4UnH74c2gB98iQLfcapzDATNN7OpAiKgqDrAj3pfmy6xZwdV99HhWS
3vlRgT1si6lOGzBV98OH+ZOzrf6uSpWao7hrAeQO8Yy/s9gnR9YJeN9oH8KpvpyK
4z4Fo7FUZ2QbB6gErPIipcOIX16b2viV5mbIHRuLzs1vr2KCUCICGP9y4Gx/1M1d
C9nbE/uzP7puub9/mmXj9A3a4IWy/hS3YYufKvRm+gULzF69Zg8FD2g6wk4QpthC
dWyvFNH6ES0Ugnog9uRs1bZm9X9GDEvZ+ECr/uzDbeCrkzfxHywK73t6xovOeeCo
FxKT1O2zMwvy/qjzTwGe7JBGmwR3r4oferhMPlmcTN8T8pcpXIOFji1+mcZTWXjM
apK8C/orGIFbJb6Qk6g7BYZQaFsg0XKvxtvMLBPOIg4L9Dcg74N+5WUo9iBhI9Q7
ONLi01QLcxLgtrw/gsuvsv144bQX3tmM7io1Vku2x8bRQPVJD8Ym7xv1iXuTjrfR
s3eICYMUIsV7wTxnnQMTham92cTeSJ0djYEhVC60SoRPfPTD8Nc5ZOQTvte5mDZR
e9O/HmVkwHkR3zyCdXhrSNjtGECR2B4b/YY+2YQTuhAJ2XzD+J3DYg+aCeYurKIK
sf4r5yfXI3gi7I1+pY4f4Br4lNV3wCL+0kViQp2B93nMex3S/RFxJqGk69An2kXo
AbZI1z5QvWIDP5YyFM5/h6pASXqoQLZKgW3LkRn3PhSsQvSn81XIuqMePDpUyzKL
tSU8TBe1Vyx3/423P3vqiLZc60VAQA07t2ZlPe7qdlYc6k3lszXeFC6Ie7zzt9FM
28+TiGgwjzxHwvVGqr/fNL06RY+SYuxCBWWdx044xyQxfttdQMMplERrpHFc1uPR
GM/vC+pyRYedLrQ++5AviIT7Ub2WmPeqm6ueJScY6fx4w+r9bMmri1OxtvEFwj36
X49MKCzDukIZCWQlnx/c2cMVlRlBPcAVSYSUcdPTi3wQ0yNCHk7zZS0Aqkf/pI9L
BmSgirLKQbhe0goLJi4zOZnP4eGBhu9W/JCQtmcv9XZ40StDZTc/vuhcXDqNoDZj
cqXU4IfMcRjevpvLJuzdxsyycLjg6Jfy7soe0VRazFWuniHk9NuNTPBDqP5pDL1l
C6pCJ/cLphYpspgDjl/QqBljZW9ME4puqDNBTxWCAipdiqpo2+1DFWAIJLOgDNJW
R8nc2XXp5Ig4yeIeAJl04Imj7WQbhuHmQeGD5WOrEAqgnF2mB6rfVafzgzx/oYL4
nbwL3cyOyUGsWEHRsS83rE6/d13iqOJYvs5er3W7Winnxup9wnezllDfkS0WIAHh
ci0yd/FbBD8ZgQUBLC5thfT220kEOsDOFfrTcLtpl3tkGPqltbmpkGUkKOR7DRak
O27/Toc11Fyqa63c8p0OhvhfeXjKsHDylu2oi2OqnRSNFeRpsIUJtvFSU58TtR8I
lfLJotOI9bS53U10Fy0c8e78d62NO7X8VuUaLGyIV3N15/CxkUHvGUjZ4vryF5hj
IqawYXxDpCMz8z8s2pdWxbzzJMOMyBXmW4pZD/CTxFly4rR+YNfkU5RXIaH163L9
r4JAHHsA9DZm0yD9RIjxhfJmyugHNIb67GMZ2qrTAIlYCS+k/nmY1d3Ykawcg9kw
dj3H9chvrm9/nvOwNkGWPp8RGmTa7r42f2JIIPjbFffUmewy5vswvWBgRW2bC7DE
DS4XCk42f5W0QUPABqIqyrpv5rAswvIHf7p/I7Kj1T9YbpQV/fljuHGjC2cbREGA
LVKysI3i8mEwe7DaM7teosbPNMZencyjebZQNF/ADR+72+yyhh5PlmxggO9hqIzQ
MrMfWkhuMTVeZ/TpHzPObcuzjkRpxPgmKhee+Hhn6eyaMZ8wy8+V8F31O9fvfMN8
vbI1cdCUpoO9/jrrsgunugLkuEMS7hrgWYVMX65JFu6M4GMskZ2IGd/IRifBd9Sl
904YZbrfp/tp+kvBbpdhyDjk7ui5tXEySKBBIzIf1j518nfVTUA2MScHl/DEssCQ
Zg0WujeaXDWYe48xeZUqUaLqHMZbPTacKls50r1TbUY53W45QIIs/50c8/Irefpp
+94YWiPuY3IIsAU1RN1ZldTy69IUJHxZeSo73ioW9sM2torS377yEXyWM8JtX+vg
jXFu6/RZEUt4/4F+dsvk7KCZrb6J3OOVCbFuRwGjV3rigE4Np5LPf092UzUfnkzA
jDlvNI8C47XIlRGmKr23nsWcpCWdc0OWCa++JZtu87qvHNxx5+gYo9yaQ6dfJmML
Uzj3iGq6XNxPDEP1F3ZDJbEWTXZxrXPRY/u/psge8wZ/TkEV5hJi39MDJXmGm2zG
PZaj2+EHD/Scp/E+B3FXQVAklF7k05336UcF/wrDgw193iFCz1QKTY7velry8NtW
VCZpFwySPbqafsachm8fjhw/MLevRUZgBEJrRReezQDNkuFWeDTF92UFF3cWvRGd
XrfzPEAffeNL3IU4NaxEBMpyAmy95U9lIqJmb9XHWEPEuc5G1HPJtIed8OLMIYxh
8thToWKPgWOvKgBFfuW/COVRDKSOnWL/DANWZj4vCovPaxpy8OZsDHQxcK1sHXR6
FBCyT70zrH7WdAxWcyxQ8pFyB+KzYDxs1za5Hc7qZohY/fR89AGcryTkJvz9xoQu
eyw+fYCUcSw8TJpKPleNr0HhJgnTRGYxMJErpGlcgR6smBVk+UdcVgT45fmaSq60
guAZ2ywN/6U8NwPItKCWvtqd3JCnnDfZskX13iE7kCuT4fvi3nbCUFGU2ZgBQLxK
2kXU7gdSD8NhUwCvLlgDXLnQApt5FKYur6gdFL7EJI3H5xBB3ZRIEyQ7zssNXVnj
Nwm8mtl7T4W63WyWdCeboifVc0/fxWqPDXdTGFMDSYa8NmLMQwhAkjdKuTop7UGc
TgmuLBEWWgh+xCTPSHa1wNRXnHCVyWweYTioRIbP1HNHOYr2dAcw9JxqOJptIcBd
V2jjQ15U3xIygWSPoCddZAfbb+h/gEP5A8gv2fj9Y/OASQwUV0pG7zFL43w7GvIF
Ufvq9wiI7a5jP0Z5Mq5hOGW+VlV6Mt0c0bfQLAgsyq+ZSFb+nt8NKujggnGeks0F
/I1Wn3PjMrY5sYc60zsS7gJLInKmU9NZC1Uod4gn0uDTrKBOPICJ/MwpsUIdmHL3
5NR6aFp0+2X4+9AyFVQSyc8hRLsSBwT/5cYBdcURNCQoYoABK+Kg4aTHIk7oJgQc
dJw98Tt3rmy2t7IEbbzNWW0CqSodF9pdqZzoGTUL0Gg3sqj6SS3ujSc5JY5taxgm
WmUjc9Oiyl6/rTLp2M1Oby+yusAxxtGFTM3xKuRGW+iBTEQtBswJPGvRVawarHk+
ojmJY43VFOOKVZfSQT647mlIk3us3rM3cAYHa9rO0cFPFfAq0Y0x1IixsOW/hUuB
XIVYSblTxBoDAaKsTCSE29mj2Vo1rzUVTSkJloXn34ucDpSYbFfrctE3zAbDGhHl
nTLRKkrx+Lv5IHMAbbYRCIz4/eF/CKFEG0j930Dr7Kpp0iFDhVmxj05C/zMkPTau
iMmN4eceX9jVRL0pf0fbGwR++C2PQ2lwDiYi9B8k7j/J9KYC/zL5bCSbcTJh7N2j
RxpUHaY3v+TwOcPqGaLnI9NBtBXcOanBsuF7yCFwKybSMM470wE70ob9fSz5iuN5
GLLeErF+9I84NNN79dVE1Qw3BruSC7s380F/nIytxpVmC1dMKb5FoYfEblrX3Ze5
JVwA2521aClzfaV53sLhNcpBQfOD43BBirisUpt7IQrtw9a0aksA4sxlUBd3P80U
zLO7clejludq4U5HLxQR2PGUuZ1PvcB/RARWc0NXAZy388PbB6I6QOiQSvtrpEPT
0M42R1NlWoLHp0YS1csg/w0UHO3+U6n9JZhBE5Ahas85/pnTi+m67QphbAuAqvAh
GXDPO9FxaRz5CHewMub5zs2No/xPTA7SH0qD2SOOFBJsYH4D3iTtfCB/7AdXI+F/
IUMeUtwtykvZLmnsK4g27/AdnCqQp/AdcFgRttb2yFE06YA0coi9uRIvjWTZi9XJ
3h/WQR637jONQFDCbrP2mQRHb3XSehvEQrQw4IvzhQ4/tWewrZsjQl99SnlQZSE/
dwjTLfB/mCJQUo6jMjmqvTF98oxMAvQMHnzVDClQapvHAcB1LfFo8Gegx1QbFYUy
ujg/2z0EXaCW01rz5lv8Sf7h31PhLBGALcUxkrbL/jT6yFlRAOQGVl1NtkjD3Gtw
+MayhQYzopSKRdTo2xfD67NiKIGMirlIgiZVMlE4+gGZgramzcR3UDhXKFV9TgQG
U/H5Ox3C92ab2THXi8A8Q0aYe2Jf6whQaWSQ/4EyAbdf5mbfRLroaZtot4Frcp7i
XoZoUdRQfIaurZiPLfbxJCiimg2nd3htGGOz9Lpa4aDK4wW9qgNqa8NGUpekH0mg
syEbJCjHJ0n/Ru5TmR/mk8S4N2RseUnUVVavl+IrscHLIRl2WH0Z2sfzSRwysJQ1
isVaWjOFPuDbVXiZxTH6s5koDSAMk3BDGMNHgNhn8KUnfAw4WrydOh4GXOiOSNr5
4/Zr+zaZsFyXZxRNUxURuAQg/Fy6kWCiP7AgDk8gvfCFzd/MIraTRJM3CGpjP5e8
We+iQBIXsctZKR6OAvfTzI85kBmpubznNFjHdpiE2a04EwIu4VboMKIwlRtyX5tl
zOpuPv2+1pxjkhSTF7uEpr5mANPATZU1Lpajz9PhaewbX22kkdG94ctRwbJN0GK9
cfaQpZl3uqrNYEOP0uq5hoi9gNWIrUoNwhk2u/ve2V9BtRYAD+cZQGI3WNOHhOHS
wr/halEGnlR0q/xV0UQP6XZ9YC3WmuRf8C6FPh3nXdPCX2vli5NGly3eU829heDv
G8hquarvjX5n6cMchAneFiL6cGvoJxEpecr82s2mvQCjYYfB0lZWD2/QXT29oj/s
kTB1IWUGBD/hR6js44bnCYGWlw/elTqXxcG5KShwZIo192lkvyw2qYMsUL5bF256
+ESMA+hAJ0EDPqNbCB3NTy861a22K+BAz4YvT5pRpVlACz46N2fPrWiekdP38bhP
S2mL+qKCw+izRlNqx1zi6TB5F+v8Eow+JzZQwLLbQ1C7usyEVqx5ivNCw814u9BP
pFwi7dXl9bRg549WYcu0pypUW14iOvTNBxvwKwZxYMl5v4NpGWUFJxjiIsAxlIb3
O4f4iTnq09VnQB++8rmme/TcPXZU6jV+37wPhvJ5RTsiLyne5AfWv7myL15Inu59
NVOIOXYrYOzyg9fpdzkS+Jt9Qjs4cMeCFl4xMuhKRwMklaBPAzGxnrqHnoNooPcp
lPRbCyin4y3KO+2slvTTIcSQcn1RDP1AQ5z6aA4tuj1CJj8t3PguMP08RUOI5KiE
rZRVnKQqDP4qHdwabN35CyoSHSZdZYOZ2+ho8Y3joBEssFnDRR8vX1XJqJCmXwiP
+E0Ig4P74vEQ7F8yIB3vRjiz8pp8szYF/BjrmUL3bMdEVgSU0dTjute/Ewg5QTji
acycpWN4ePdlgGNujNUc0clpnzV9DM3k14SHadDAj4utKqkM/WWsfR0/GiPLIlWj
sMPx2gbgUcoPolvxunYdqkb/l3davFtIpBmVsOs5hMYMQAI3AP2tGQPmg1JFBkc1
gcfjbYpFQ2jVPP+nqZqASBDK5V5pKAEuQa+v2nvSwMRDOqBEYxabi7XygszfVUsQ
zj7yF4/dd9lMn9/EI3FfJF8wGIKLP7pSzK7rhZnE1uO/1rm7cTWpY+kYNhEJKY02
CD6fzj206Y56SzpYkRqUyI9MoNxK6ZOzSe+K/LxGpKvxzJv/fiEMnt7J6n7pCCcT
9pRASX6S8V+nymYUTXZKlT/ejgAI9NtNB41uwbRr5zwWEno4PpvmI1qTxGzVBby/
ukjtnwxzOF+hNhPkqQUIG3YRNJX1chlp+4QVWVSflxfrfIsEhc5fUQ/iVolp2mNh
EnxWH2HgA8toDvWJKXPRsdPWs25C6noNySAh9/TMCum4dkQyBNnnCY7riOylAmq+
W40vc+FewycpKUfPm9Aw+ckbBYUBOZ8qyHGU8VKe0BAmZiXcvT4/bNZJ8Px/r+Gn
vaR1AddZdxXputhFTck7Of1SNpYgLMzMjYta17FUv1iopsRUZuE2FNEvNIKTrfCB
1BbSjuNBJvsgijaxcQvhKNs27QTZ9ycoh9RTOqApqK51s3yGh1yIn/0I5Fh2izNn
swDCyWM68XktILCennhzjG8/PZTgNsoJm2KfYeVRdK6gVRLskeL+c1O3Y5ou7RCd
rmxVzjK8M05MbPrRde8IkOtNtOPzw/+TRQvXk33Y0pfHEFvj7Iie8sSWK3eHVc7X
UllfTzsax9CHETscZwaX0kKYUkHqnbzITse04qAxfCu0aopnR/z4TKfgponc+kOC
6qn/NL43TuZvmaRUCYXApUNhWMF6c+Vkr7ZhH0ptvUDq5cRCL6gqzuP/QFAfQJqc
nppdTenzAPsPtSypPaftZRgOt20b9TovqDXwyJSd5QJgA+r1fFkx2xsXXfnasEsV
imDkhdz6jpPfMq5tR7705NQbkrXttCjGelwz9Mc7Sux0u19LW08a1oIsL37VOMfW
9fER+mTFS6ugPgQJbn4157oww589BFZGwsIE7OvgOuTl2JDqfNnCXwDxEsqdnAoh
mTMhpKz2xwCO0mYVq6+eY+gd4zPo0pLyB5hm8ThZRHsQinrb+Xyf1NkJlzK7rsQZ
A1H4k5HyMjEAEpTOKaFyDeb8UODRsCjIN316VR1d0WaycrzadHvz+9jwSjX1ldYu
GiqZxaJ6iWGjp1V5h4V0HCJNWTzswlkkHf1qrrWlEBDbPRcbAQtzYIUpd/sPTsUG
LqLvW/FlQYZopS8ccEm9mTLqqIRttHYsoqGfbxGEuoHfAtcVqIg0zF1kTGDBMTx/
gKUeOa7IIAPHnP2EjvDSzqwCaZI32S+XTjjscvPwsEQMItkB7us9BtGS6F6adxP7
tJGTlETtQ5xkJQtTLLvvz4wzB3nQzXwoegSSa3EcZpamEpzvtfrSxjLakwDYsTZc
xjfoerDwhbBztVY6P60Eg02w3zkkggzA1nG8yLykUou9Z3/rMiN96juMvxsJPGPu
socwB95ruRvy9DLQDq5k4ibmYolEsObL/ZYXfTe2njFP0M0YiE2WXl5nLg5gpKjZ
oRYpUFYDp9ZAAJwxsA7UOAUtrspvjomm3XigiUfrFBMkuwLo28lnFkzrpIHR08Im
389THtVuDC1VARnmIT7l0f/E0v5o4M91b3hcYk7u/YRL+ALua+g6ZC1LpAWmzEA6
XyLB2QtMKyHyHlC4UTkVfGKJmigGvQIb4lJk1Fci8yFqkwcZ90vKrxMqeWAsCOW/
a2XgE3GNSMhU3YEETZrpmBuig1niR/9jpC7w4PDrGwpkUpTeRKi8ic+omd1l7wVL
2Q9P3emOMqCNmKW6IAf1fxZZOQGTrnukNMYprdviSTSBuEotzKJQ3pdZKmM4VKLm
F1Tmmdod7nv503eYL2iwegy+HHYwkbRKuovdddLcWUu6l902fxQxlLnMeFn4VKpf
SR3HQpoJBJFm1Ao3pG8drqCktPlCoOSnBT5QvyLG2561D1YWudjABc3CO+Io0Tdq
r+O3Rg12G+uZc1lohlxyFaGAjKc9RIKQZcUHAX0lmmgI4OshQ1uNX6EC+b8hqNLV
R9u7kPvXCQ+y6hJo2z1mfax5mmyISRbxk4qrljdLgAbKM6p2luBD8Cac1JvDfv8Q
Db8nnsFwIk4rwfr7JkD7u0uJTjbZTCAxHKckB7DtJXt+foadGfisujmdOWPfzQrX
bbcxNysG0VgtuBwHOtvF7YjwZBu4vUvzkBO6wgPisqlUez7v/mQTEzactWJvX3/W
t+6YX4uTiOLU2lhAssCBdVL0Z7qrV8lvFoTKDfk5DZ/NUmEE9r7esGKq9bRxaeJj
3LuBZ+7thPsfgp0Xs8fzpVnCFy8oa0ZFfbyMf+f4vIkRwh7rUcoqDKtA35i1u15K
yKaW08iBVpEk8vnqZQTx9vtPaS7CtlfgbXpXaiT1jsHxhPRTnrtMB+QXdq/4+C8C
embiidg13CZdWXO6Eu3PgKyQKGs2kITjST/FHZJByYycvE/rGxauzWEmm4soqBK4
qBWeICHt1wA3iocA+pUUiiqOM20DRQbCCJwLoIH8YOdhnWeuXKWACjrA0wxPbblZ
7Lb2aGGxK4Ici9h+Bo65Jj0IeLttMpQPiRfVIQemLJYzjNJbrJISYka0/zfTXJX5
M0ADFoCnoLEnXVKOlFoEKZ7YQy6bTyPOxkRHbKmW/9m4bOoMyP30MNj4P5lZApOd
uAIGITe4J1cMzJlaTi36l95jTCT7hYtise5e03DkfpktDtbRNRdpfh31+vQ76Eff
gRL9pQtDY7+B9YHt6xcJ5HgRmoRomctA/gbNXOyYL4GWhOBAlmxmNDUhjcFIIKZF
zxSvSn8QGfOd+LbopKUx8Hzcr+7+uzo6+uRdSN4Z3ow2v9bgOhWvXeO1P76x1O/p
D9GknYTCZjap/RqmluRAwUp5Nq2IPUzebg+GCtCi2ksyuLmwg/bIFWU8a55U6idt
UGulvivdvkUMN63mxZXqoEM55LkPY5zE3OhxudcIHLfnogPAwAAFMmWx+hbAGHH4
fXuoQhdta1dXg5cPjRPXiSD5L/Nt+UOdT85EmndNBLmiUDD88vnGJc4zCloeFQKm
26KdVLH0fwvJ+vxkTnTWS9BIwQlj04+NZ43QnmTzd76FNO0LBq7fIabE/TEqz+ni
Y2ZQbFYAggWqxKi4z8/dSW/CLYYuY4g6ktUZbiZ5Za7Y3S3ouYQwOYqzVJcFZ5sx
XCqBsBNx/ykx0XRzZ3zgQxmpRiuW/ZOfW09N1AOSuZQmrmjc8CIdijmkkZMQxUrP
gzqRA5uGyl85n1QP7DGxto+CB66NIBrYXAdND34xkUUwmLF88wtQtXODk0DOlKL0
MFgC5hnMvpv4olibifE0XiCiad3lem/eCud4kJ3u1/liL0Gb2t5I/0RLfII4wTPr
t4JkunYTEiU2k9nkOZT26VN0/uQChy2XY1V5zFOSA3V/usJp4g2jtH3e0IrTsKLt
m7PWu0nkxGQUvSzqsTN9c9tLMimAG2W9GmanWilP/NgwEvdSztAjJH6DO9Jy6eEk
HnT9aBwZ/dzMGooEdfj65HPktFU8wbp6a7DwjpHmHSFtZHblO5/tzRbthRnd1vdE
hXscWl0sRJiwiKKB0bIPjY8OvvhIndU0dnMkhZtot0FxtynnWACjoI5sbgujxlvx
60UeskdjbkAg1MbKJlmDmXfAdAXTdH10v09Ujg155Wh8fxh3jJmJh5aRZ5OR2aJX
91DLyV2W+px7gIWz/PwZQOJrAAws7GIfcYKMraM5UVWORvOZ4u6E1nJYs+TSHOGm
25DXUQk5laGNtz1nBo0GssXbxzzEdKqAViIOvxSeNSinYedW7psnVY7Oj9b0KSKY
kdBbSj1JYbOoI/jTw4dK1EMKU1mt3COgxoIlMOrmTbOuhg+v2/K6dueR+KLVu+YM
snkDR8E3qMlSAzW94uO5bzHQnEAwMGPSLABbC7Qi4907aCAv4AU6f3WX2bEgwJFv
nA/1wFKLKXDsZlDcdpSTKIi2/tdwWbl6oV18meGYXnEyFACMtFiUAJ86rKWg8eYK
62yWdMSJB6p9LwImj4uADYsfD4tOfnSEQnMxd8FryLU4KHledN+cTJmq+cuxH97+
vRAfONeiXA04RkN1dH1+f/aIq8X6up1a00zU00GbOWbOgJSOZe3xuVMaf80wSXJM
jIOC8wPlgSMitc/A+2qGvn6Me8FhVHEjs0tXulGV2FWWBlmLOI7aWvmGndJyBB52
/S8Z2/035CgXFyNsKFtohrONdSjY1mfv9M+grp59i0edyZr8Y+QbhJrI0j3fmr3S
8q01U/cqfvAtc8q06ALldoVeUBC0olqZe94M9N60BPo3fd0N3/LsSp/RVz3yrPPe
QEZ/dTwctdLDFiiJTxjfsU9YBSO/m6oSWEVkBOJsC+XAB3XSf1bs3rRL9HYW6RXw
aLStSxjp/LeIEYRIb/aJEcoIc0vY3fZmqvdKldxBebtYhnQrDDnj5WuzcMR1JjG4
3hdgVxGpGFRUGnCwiWTo1yX7A8hOLCZFjilkPNq5jjAJL2hHnBUTsIgdfTLlMWyj
4nWk+VueJsFNlZMkhynBstTtz8ceEeeKKelqop1tEK3RAV4YmuVCncMGXtK3PoMn
0Iq75Rv9Oof0FrmNLXwgUS+hLlIQUvS/k6yX2KVme09miR084/zlyGI9+D0pO8/Z
XKYJHSYtUQpEirBaaQzef2a6v7PYfYoy4H4cIN8/wrvWvKu7rQJE9yevZm7/nnef
C/Uh7PFZz2e1nAHgeFYytg0TkgUQidOhqhcGPO2/HeNTYVkk4Reb0PkonlaTw/Bb
XvUvkx4RTNf8Tw9gfwodZTSwIiRZsPNsKrZj716d3s9ZBVRaYz7Z0vt/rC8HijUn
ahLgxhZduVEKZ0uMW8dZTCjsipvoyNdcEbqO6UvVDRWZgsrF7tSEp9xw+YwyTj1g
W8n+kD1RrdC6zhiqpY178c3YDxL4qx0R3GJ8uxYaifkZg7vt31CD/aXzfvcTZfl7
/tSKFqB9qqjsr2a/UxyLnE9cmSeXHIWFNavdLZNDIqaulbACauFgUkyiC29shf3X
7LigmpGc14pm43YEUWwtBLgZotMo0cxSlE9K0jIl5fdnjyLuW39ai+r8C37hp61P
WkwISLz4u2MmZfJsvS+z6m0y0poDa9gIxF9irtEDjBiJqFvZh6Rc5vaaMiF15jqW
/Yhn3AZfDVCRCxNzkd4FowMeK7GIFZkP631C+qFSD9zRYQgmJ5KK5qG0df/TnPRl
bxIeKJjpBvtMYdlVWmm7Vt1xDMl4TCR3PiA5U6OXcQ5rOJWQ9oe/wztjQs9uUfPb
27Pnu73R3ChzIRKqKRpZGZDirBopBYrTOY/8XE36NWmrRKKazwZaFpEjQdTVGzc5
Dv9lRGY/HSfoVxbuSRIb7SzAgphJ2IoQa+nIo1/raS71y6cKAsdV7ubP6dkOnzP3
dO5sAsaR0rMf3LelzDVhvk1DQsrqrVhorr688jK3Cc9tgOZY2U7252c9f5M1TWuM
DvGcMenESD5Z2OfEhmX5A04zGW4nfSg4+Fg/A7lHjIWfsITKHbUqe87P0HOqR6lg
hchAKS2ezJYVcmcaLY/6QeijAN3TKZhDGh4JiUlZVq6IYm3FtB7y41MWWf/8vLAB
OWRdf/3e+3JfKl0qN747wP2QDTSUSCkGciVr4LAtDRTPn8Ig1VQR6E1i5BiJW1Lz
IvjL1hgCqlQomzrcs2ROnamHchu5hiSyo1Z80pDsH9fVhArn/SQTnOlNjCxh3dHZ
wFZR+mObK290c0IPfjq22gkO9HyVAxXEZDSLi4BNNkheYclLfO5toBJ/EsCS1r2E
SuvoqzBrFKTMXMW/zw5rvKddjdWsg7YLTKL+TF9myW4onFzpVvMOJaAkIf4BQ5A3
Ac8aVXc7ZX89mbB3wQGRI76HCGFflWCgKUNRhaEuEDPp2BJtvOJjIEpUxEHzaz8r
sSAxXmrsxJ5diytyf/x80VKmNcR0pLfnSonX7ztNvGgtYnsw/kuqEym9ffhiGzKi
Z5t8dPaKaqPxzb+O22w7PDqr+wgTff8FrbCUPbLLeRyXbxUmke8ZF1CWANBfsMmi
S2DmQrMZyA3WMrCMtdqeUy4dVkVFWsVU1sI3Qf7wAcrTrL/+tzPqR3I568VYjwW4
L+gdXDRMZ7EafKhq5fRkK68b90sPcB7RqT9A4j0vhvL+k1K43uApRGuQYSFX3NU8
lUN3KkRwpjE66Y7koXIiepiL6qIkq4ohA21fKuZ2aD7SXCrdHuEfe4xPwA6RcUwI
vFWVpBy2li1ySYOCYHijtM5/PAOBs4BHgS8WBa1KsCg/h8BcxK1EOmCX0jXox+DJ
xN4MfLDYlgEbCTwgK4ASiBmXd6Otp/8ZWZSx4DUcYgiDcAr4iroiJiDt4BjXmEM1
4SxEzJaOiY/Mc3ufgbSBX7ZcU+/kJPaOXRu4EStGts1BrMOpCc83leqCmXLC7iFa
E+iZcpBZoNZUNWcS1RA1vqzhacMgdHB5eeuG9bOWLMeMim6q02l5WGChGUVebgz1
QlyHC9G92lYNe2JZ4eGTpl7IYhwhzghdzihZEjH0RRGI0BNVBtfgbjnnvCA87DFH
j2POE6VWrsCuEL85cvn0zTawWyR8Ue4xGZ9faP9i5J3+Ksb003Za45OG6MvUnFG+
S/t1C7dIHOJPEoUoWrtG1t+yX3t9D1vcpGqPT8nKRqlZLixKy4o5SYLKYB3mHD0v
t5uvZ/xMp9L5kTNPB3gOWcAH3vBXT3JVKDQCSRShVnu+rRrDBKYVpgsrR0RoSS6j
H/Yy0d0DG4S18Gf4icSr5RCsR7nxkjj9QX5rbfyokgwmNL+NyfEbZ3c+bk/TGFp9
ixqBDITcyApwFvy+T6PlGo+aMR6Jo47VMpedQ4gmBVYkq4JdUKJg6pNKytwz1FGV
uEL1RCzNdI3SYtuTJuPpsjLOUWfyLGkedMlsv8+Vv97yyCNxhSu94vYi4T9f+Lxu
x81MsCkPNh5uIHJmffz3OEu+YhK21zTBn60kzsdbJ5QgVpEqcsxXBv8fesvxNGdj
b4fgD+Rdf0BZDG7CqTAs4HMYNqQuS4ZLKulVk2R0ZmULVx7x8nBeFaEr6QUcdhRS
iydiiVOnUHRSEmk5E5nYGUo6c67Fr4h88Uscs7llB+c3teEfEil01NfMszh3ZajV
pOCD3x7R5/9TyMHBaGYfLs/7rAr3Js2IB6jjPFtq94UtSIDTIirtcBd+wBRNQPWD
e7YswXjVYX55LVjUnIT++P4lEgUzgTyPDXk+sbjfWllUwVtcI9DziVv8OZ65uaUd
NuZ3wuOlpLvWpqdpAPfLdbKQAcUXnr6pcpYyIfA7U6wAyOizBKatfoaRr+MJTx3O
ksjk879jnIlAhTY7/7/+Na0WP586+XrZw/XgIJn7fG6eStLWuZv6zDQXfQji8uJH
EeT/f/YD0QLNpTCDp+pTwkDUTmaYtKeMcdzG59HmIrtPkLhLMyRu8XVBDx1oXxiU
7RkYkzBeBBbzWrPS6lnB6ahXQ1+jnMoIn40du/lY4CeziHynmghmtHsGq5HejElH
jPN6p1Pu2+XpnyreYEy2wXxSic/cXrabLEfXch/zHApLoF9v81fKFBss9N2AtTx8
V/QJZ5TfcU/AtJCxDQ6FP4TNHQo9mZKrsK4g6Lx4m+sCmOEtDfPH4tiCw7OxuH1d
2CEGB0FcmEdn2OzeRyZhdjv0tW+c8zyOAaR5AUuMSYesk58bI0212Jzxff5OwqyF
bYWRiT94QuMXGVKzoLWUsAtEp759nm3qEYldpUxWhtiVP4oxHW+Z8uIRVimuJ8gy
UZOIZan2g8saZdAj8J9PKNmarNab7bGVv+luzlesCN1IZk76hofHTeKkhCsK/aaG
vVW2Yw9Ryi0xgarPghMnUs2rLknzqpB2D0Fg09johFQUw/ODAtHi2YhD7+YidFgc
tBKLal8fWIo8clXl+I+RHGJ20Bn+xUwL14HF/vmsKKSWMoMFcq/sCtmQysvuf6UK
oJWh+KhBxDiS1G7scqSmxECjKkhEGL2FH4sA9EeNGLDoAfdDKzrhgXUhmy4Jktdk
pEsTkJv01bubQFERkCoTtuPPht0dWfXCJPDOyW21IHSxPmNyYjhzHO81agbePOtm
YPClStRmlcXr+iEkJN7liBag4HSTndBJakr5Rxw3EjPHKPb7Ev3tYVR5siumoonu
buaHk+hR+xessco1SOnt576htNF77XS6OOJ+YLp4SlWRRAERzQc58DniK9BktLDs
/t2VcX81U7aZb8oLbGXQ2xIe95ZGnEi2y9JKivP+IbqFa9tip8W3C9bw/+zjYwd7
4gUuXH+cX3cCOWLdG/rkSss3GidAiiqn8OY0YnJ2sNazUXPg06Su3zLL1SgEn9tH
9ExJxgbCS5Fd5MbtCKmdV1yffCIkj8+xuvuXwkIxiby/PY/p11t22r5uw5W0RYRU
/heOp8Zf3dEkUNUXAIh3JiKifT0NHHEargNxIkovcYMBVqybkeoLkcxi9sNVaOQ5
cGie16FKWjGMYpUP+dEyUYc+36Kyb5ezfUHuWaAkoesFUxzYt+S4R20sQGPuHtCy
jcm15yhLYW0B4wcicsc7LXSym8EuIe9+SETx1jZpv/n6x7KMAvwKcusDGzBGHswO
eyaDZvyTZ7UlSOFhhlS+V+31IAIR6fpf6NrWOnzxcxfN5XI+ovLoXSQQZOgIGYbX
m4tJ0fo/pu+K4OsyBBowlWpNhOyNqKYaxy6rFsVo2uMN9mFVca9uA1qvCLY+O8EW
8GxRRpe6fBLXn/KDupTn7nke7MKCqDVKmW2PjK1NKjfefntTqognUn6ZBDB1hyPX
FoZcoJWJw+AVwclOAp9WM/PY9Fpzx3zbYf2ar/mtOlE+vDeRz5idVHTZJ637pOAv
NpNPfH788CqFsGMVdsRbsFlzs9xj0U6qKxdwdU5sMPDxSZxLWPlx27E3FLJVFaYx
gZtZdG6OqH0vQr2uJFzfSdr9Eoaa2rb0XbSFQKee/4M9UuGXkh3wZla+QKn7V8mj
+yLY2YnqBCw83IMS62DHihZE+IYllAhfYM1NXQdmLsFOSxKx9sIdKkhXUNCBs0B6
tm+Slageisb73fLxlhFFN4hWbkEY3cSk0ribvDqcbv0FzC24myH4FuvkkyAdng1h
6uLSd8JR8y4bPkjTxkQRmUQfj90ojLXzz0JXIc7t7SvPb69yuuRGh33qhanQSles
axWzelZiTlSOXIPQMZgwYowQLgmCMQC1+jJQhXoxR9ymfPyO3BpFAfHfLqUGYIzf
Vl+qbFgOPoC85ijks8nJ6F/kec+UhRP8e1tz14furRwPtAd3n7a3XhZZ8t23bgYB
sz4HBkxr1wEklqqQunXqsB1hiufY6PmePGElqQnaFi5h/P2yUUc3EC0brdY9AWhg
d+B/nMbrXT6XSOZZhdetf18b1uicbpKz5DztnLjli6BS2eMhXfiViaRdt4hXvjht
H9derdowZeJtsCQ+ykb91E9r65XpP6wWEx1GimivcK7MODHp5POLs49uYZjSKWt1
TSlF4qfAsabBji8jziabw4eg7f0X/iPW1cJPCUQSsNBLJaepqVJ0mUIIkumZ5mo8
pToNcvrT4nrSTSjxQGe8TdOxqLDLb3tUpqVVgCSB3Q/7CU+BkyLePCfdf8f4kpD/
lgDToD+F48n0sL74D35AsdNJhiSBZhLVrWG7O9tlarQ711L0MFm/tQ59t1yFBxlZ
MclWp8lnKaYhXBgFc6FBm4w/sF5SohY7ZSwPKX7dJEH23ujtthmAdSF0W1LS+PMw
0WOAEgKoGOoFMJ2/qTYDJ4kSsamTXZdtpjuBsYd4DnIEwZIjQ3e/YxtzfR3mzmEi
XRSYyfNfedlkyyDZENYb+/XYgKSITn7VqMzCTn2mtTJ8+GJ4uHOTNq2jLw3wGW8A
W/X8xyFyCkoMGXu1u3Xwmv5D9F5WxR8KGNqIndIc5LfSMw+dfStxF5sl21Jdq+O5
+uucJui4r6PDRCeb/LO2ukE0nFh7IYFwXAv3spozyodW4a/rwNmDSZV6c0O22SBg
j+fjDqmcWbcjuel0h2yelvQ3DxyG3ZMWh3QV4LfR8pa31eHu62KXsdahFVXT+SGq
pvDfQgqJMlAe5QyaBQiNcmvGZacPemTE9AI4jvQ/nVHLCrBVEflg0TYJWCce+9uZ
jdeCh+ZVGnPXaLxTEbNlWu3S2pVIfpkcka5H3aEq9BydzulbxJrWjtS6YPanPxo3
NfHfv01QHMgkpphUWtnuG/wlgACKjFlohh4s1MP0GO9nqaI5si18OjYXG0ho2Eke
SlZ5w9SxLI51UD/tvMOqZNjgQdBfr3WwGJJuRTByqgIreB3S14qknSrZnwJSArl6
7/bxA7YR+bFVgHmPq+WD4rBbwsOtgSyDaTEytUte750YKuc06e2o72ZnceQejyqz
X62l8OkKFbKVGlGBzJsDZHTTbj9dQ+ZV2kypE62KwCBUl++8NOUIaDf/XJkHexiY
QalXLO+Fr94E211KjA7K+7D1bniDSkT0Js2du7QOj8qtKEmVedEuKaYiZHouIqLZ
AqstaW3lOD343vejGd+3oUg40c6Lesa7CZVUzyr5Ire2+p663W/oU6b2UYAOS5Ao
5bo/jVaRPMyt8UBVqnSl7tW7CwmWejbtLU0fyGzoQE53Vh3M+zxJ9jxl96f29ccs
9sO9Y5Y1md8wcT81aPSWtdxIoFIdBJFPS+m0DESPBwt3u1ft3ERJvH3Nps89pVVd
xOiCIv0dmizPWXWlpqbu1CiXC9GOyf7AjaPicsLkTpnaioqYEOa6Jl30yHq9xfhb
uG7uTAPQHG4rjbBJgVviNTXWuGyT58hhdG+OEuVlsB/0GMRh6tFrZGDGSkBABJkX
GJhm/tqbNyCGApmWG8RFLtna5Dat+ug8OORt3ADsZzeizW9EQmxTh/FXZLZNx7MQ
wmOV+O+RmYTQd5W9/DKjU3F7K0lv3CsOyPs4XPgsqK+wxndLjZM018eBM3eAmnB0
jxy4DW2bBK0Aahrzd5Onb65pHts51T/YTCPy+5ocOKJ5DJbCm0a5Bei4aP5nHJEx
XnvgovTy0gY5qvEDhDX3P2g4ZYCm/bFvrLEJSYOVla69MyOHr4jglybuC1MGgwB2
2uMQ7wHEDgNdINgTwWX/ufAUebQ1hJVjOdKzt2aezgq78Loj5K5TFzqgZNwyQkvh
kDwRqQqjsgEmCmu3LvqyZ+2wdmQo6TP2YFX6eqF0mLfkNSvJZyLoj4ZXizrtSFAO
zULWu6VkaJ/UYOn/3IU+T1VvRtS9kJQQxkNpt4GHkMgPln7wTvDnJZIRWH4zkdZf
JGgTs2ohujroP4LgKkecyi/n1epH4Xz5+3wwdhJzUDQggubay5DHZCPXCKtW2NlY
BxDNJPEoXjfLIyVSZBkkikspKGKpBrF+q86Cpi8Db7geTDljb2t35ZzOMLHBWgHX
tYDcI/dr9lhux50h1RHAi0MH5ZBHQTHHd2eckaN/3615w+IB4UxTSGVxM1wqakZL
q6wCxg+JjqvPak6iMh6iFEsU0K//R7uHUUEaBqj72WZb4H92OssgMWQuWDFhItgV
jPsVS6y9YSu0qxL+s1bB/b3lEh33ptM2DA4jKZhFZaDDX42bwX/e27PDRLwbiA9l
lCyemee6EdmXzT5vVcQeQ2CcaoHtyOAG3hCV6JhCq9q9tFHHJNY5LrNeFJ5mSGfh
isEPQTKBVCZ4A4fe2nMJ6QGnog2mkSRtHlQh8PMXH/vn3EBPOjOjfZCmy0YiUDFb
aS+zf3goC38U92L8yBRtdwkliKQj3qTgvFac6aME8Ly4EuPcyLvYAJ81tZHjOaRE
LIz/Y3I4PgtydJkqpHFOhpAL2WXvuv9JHUnPctRWdbHcwvjIXIowvAnlUNHnTllU
jV6edBvmKr7hL2WcHaikaZPNgYYM9wcqu0gfIFE6r6BeifE6vXPKI6GhcyxK2/PI
cU/qz0QD1vKegmZImqBTj8OZ4uasDQ7Iqh4e+77Sw0/A/9leKff/K0dDhj45klwl
LrY4pByescGL51w8mo/c9/U4YYDNSj3VtKtqb2/tyNeuiSZacjrHwFyxHOFq3oze
12tp0s5O8rmL21FkBdfioIoXPSeBTrzjO2dHAp2ypt6ZZ2lWGE4wP2X7iVNLPW6a
bZM7T1wF/3PFA94Wcfs3nHjpIy4UU0nu7BLPkFFPIneJz+Mhei5E1nvmWgdVPscn
xkAkyyev8IAR4XIEIEAi3pt41aqvzOcl8614UaARn0cMiPF9JOeKXT5TifmSttII
/tYNpwo/YfhiBtvlDulSrVB8/XkNoHJxEV1d4daZ5jiKN5gUtPIoeQi/1wy8m9jM
7ROHapPOXNBsV/BgKAzPliY2w+c/yutHsidAfQY9/hCVe+oPV3Ey4K0RZdIpu6MT
Wd6rfZ98Z0wtTv59REc3zQhaqatA0jkDQ9mL1BaptqrAe47WfpYl+r/BDiduo8Iw
9ioSMgePTZTWWgWSpnxwjPGcatj2xrhm29sX6/d1N96vYs21lE3YxqVjoT6t+0Ny
cSUc9uI2oCJh1xVMoy6oR7ysss9Rm+oTO2NTdnUBqTs8nleELXDz854UHiDCuaqa
9rFPQq5KsAnicDDgSeANVbse3dv+yXDVkz75dR5NYER/gVT/9BJ4ibgeF1OKOFuI
NcrroB/Li5d7ZGqneheIyaQTMtmdE1jPmaUR7fmTUAof80jdpH3e5SQKeX7KucKz
GxJns3ijPB8hOxxMJx66HHjqrmF8YfxaEvk1rVtpezvuJeyB0V3qI6TKwUuZZfVj
jI/QVv+KYKDpNQrmz+jQOq0nYjlWg/GmMFJPUVB5a10DkoQ16HzpJmREoY1CubNE
7UuOLlOwSbFKQjZRICluuxuPnSpmiVXNc/y0hNugyIv3XNnnEWXCD7z6G/xy1cdU
mb8aZ3gXTGSgrTr2MqQ37iuchmNIl8Bqz4ZRCPPPAy8Lj+vnONVv2T5NHIHQhoKL
r5JXlR7cMA21FTmdMgh4r4vnekOCmE6fVJOHykhIkFwyr50zBTTw1Q/EwkItruiA
LobjcTtnwNPe2t/LLSIShaRT/vBWqqHm7eLQ4yfgg975ifbJpKzTggbHCjkCo2Cb
3Ax/y2RmysdqlZ/xNrJ4m+eDgNA073fATbg1bTEeHyv7p5LZAM+zH1GfpQuX5PIm
7SLE9QAnaV4TI4yJ29V6g4vSNcxwwLPTf3Lnl7narejZQMeUgWEyBcAV6TSPHWYq
cYsUumF2Cq8hiOciQ6J+SZU9mMIK/sAIKKLLQZDte4X39adXpmskVs7sIfF/CYWV
5ndf9gDOL5JEHzHrl7a4SWZbouaQ0yXfSmDfsz4FBUyZLaWxKmLw2BVJ2z5OiA3U
9UDUZDgbIMHprRjNZNeweRURivp/KLtBzBFsE0eCUNF8nfzouOTX76XG3G/v533O
U7pVh8P8BUJirGcTMyiFisulQe2a7mjuaE/tnNmgBTCK7ZcCiPfBD8PvWNDe9Mx9
RjSk6OamjrGGukV0XRx219PYXtTxToeszPIORpNNXh5HoqPK/B0n5YrZdN3iYwGZ
H19ypbGcwBkYFV6NVQY0tGFQDX1gCtMOX5YjZWuClSUGQDm8fsy7SNOb7vK0+Uwx
FsMUUxY0nCG2bLInDloSX+b7o70zGEOS4I5C57aiWQjspC3O4gNuF7UObVbWDDb/
fJ7syXop3j6ibqg9E1C5VTXBCKiwzRjUyl2Z1MnBBZ3AAf6ZEqw8y1Al3I3g5AS8
0glWkkXDYDVw+WCjE8oRvRCiK5v4pYtnW06YSPktuEK9pxAl8I4V2gwDgClilKhC
HqeQBpBsvZdOkqwqpgQNxKP4/NxwC2vDPFCZXuiNabztCRAtX8fmRWCoM/xp2Ro3
MOPBeZBkLStgqnUGN9/jybRgBLFgDXXSRMbGy+MQzYKlLJpl+rXzNH0q5tAX6P+M
6EBatDAhtvIsnc+hk/HXOImXpst/V6Ovqk8Eg7h8KAGagMRsPTuwcuzSOSFUv9gs
tHXQER94dY4Rrl6OEQgbevvlkROc47HarcmjfTbtbEtf6RIzmlWQH8ZYeFHCav2J
luiENkfWhVJgDc4zgiXDm9cbsEM2pByLwNcwxgai3H8ry1bsYWI3J81kQm1+bqeE
tO8zUD6acONN3kuusYhKQQBDWAfwVmy6E89edZNYcfxT1lF8c9M25kAecRh6GhBG
MfH94ad+zGWCDuo/a3crEb9LHpdeVQpB7EvnhYVWVMFgyQebjOa0DKAp/2JypZMl
/Bjr1MTagWSj6qyyDP7w+7yMd7b3ADxAv1iGCMerkzbHMrMunZLZaf5dy4BNV4Id
YUX2axGftaKoUlOy3nhVn65hl4tLc9qtOgA3d4IM7Um3VhPNbvRTaNpkuXVN6tO2
G1mJUjK1ppQC/00iUJpp69wpe9ZUDIRe523nEWoUghRnPAlhBpB7543ayDzfBiR6
vawlSzX4VJMD7/hdc2d+Fk5LY7Bal+qFWktQyQJZvLGXcO2cXFm0ETzBbfcCkCCS
Ar+lu7h6tg7SdbtEaBdtjR4nXjsIEHfAQ36nH4qegCfBEvAu0HkTEwJVwLoX5L73
QN0YJjd42T2qtVDFIOwHn5G6UfM3KQZu0Ycjt/H4dsajNtQX4CfQhLVmRPhV5Stl
ud/XFK0g5eIg4PMwuyv8Aidt+xhZJ1X98hnuIVsXYSiCHios+wYj3bbAm48bpDYs
06ERFXzSiAGVjsg2IuOd2ZYmAbnKtlKRvHUpi3jpzpv8PnMEXJn5jWTTPZk6JqoH
wLtl8GJqgJzLUMDYEDA/52NVzX9yvGeq+BcuRaRfupn18WixOABDLr+Et08pdx8l
cJkKudQRPepSeUlSlNPP8/K8kUekb9wrHhgdpYf1sCVrpCT/eyrbiy3OyrGKmSIw
5EPdkfNtGTxiVwdLGjqWJRAE8aSJv8p2obvY9FTlVjUEl8hutYSDQhV6rkKw8MNR
5r7VwGPgbEIvkvWK18odEJpbK3kD3n+HeN0wxJkuvqacLyLNZCjMaeoeWc0Ax4av
/p12DRnFjZ2lhCuUoYdEJMVGw91IBv8lX0ECKPQANSnuYdQa8y5g8xEjmYsMcmrK
Q0q/Ac1DT4BW0AK2yMs3exaxRGX0e7YVAWMnAR43AtWZ6NJt/YFlXlIuNucRI7wz
7DszHHnq5kZ1O95diIGx8SmGCH6Z7lzeaFuJ5TQlBTkb2K+MolT+HKrHRZC7mEDN
wmJb4NVdkTFCciEX1zdj54/bYHeN6NrQhUENwx/FmCrQ3piUAipLXkgt58cqIhHO
rMA3TNvSSWzOECeIsjN0JqSKiG7klSrZZlNGGwNVlZtixn4WbFCPxWq7iMKj44Cx
q7wuW4I/yLAyxdBjsEln8kJyL//1tnna9PfaPQ6ZyU5KsSnYyq9q8S1A292sYB7R
lJqAoJHbvJULTzhzdlQnF1Gc6c04ZQRZ17lGWoTVqe+zg8BjRC+9yNhKpH/kxPO2
R30GCuxr235UZ64e84CwoFoTB5dJCQs+ozNqGei5Xac+1pz34MxcBhmm4IoaMFGn
EdBmY8tEpLYUDWVTe9watGFmJonhQVS5DHcvOh9IkaGcETrzlTyeoumb+c1gPoGU
oqHOn0ptpfGT9HAKHcdIXXRXJt4q02bgmXkawpycypveqMtL670771uwphLSkTmH
us69yzlH+uDsGCEO7YcD2817YKuKcxqL5Qzn2u2+bp9wa1X3BJ3QhaGu3v8t5uRG
vw1PFxEAH6O3jL69Lt8R63mDAsa4v1Gp8l6WCi0rKMvaFBFhIIO/tGSdBdQBAjdC
qd0/I4bLO0Mw8qMNTzzDoF+NrTO0xkOZeunnPdVkyCHXU+DkH8F0+XIH0MQHmwoE
jjL+nJBN9+CMkQNkwnO4TyafBjlnbAVUEQK8A8RJDEGMFDShZqdlGsbV2cdRzhlF
iz8Z07crR1v2BaerVYFMzUQXZWSVU19koGSpRLR/zqFHSwin/VR4A04qTpwXyBj1
f3LRuVaTFQc/s9bp31NmrVK8SJp40+xa8JVsHhXs+ZGvx2jxd4E3CoJVsIVYOjCl
ioS9PLvfPWY9vWPT4wsik7O0WGzSnIkyj3CgwRdHe8yXRyorr2IhTcVSFOCDTlsG
QxKWgTt1ltBaOW1ncGx2ScvhS2qisuKtTLhCdjZSmI0vYIIXG9yYCiRQV7gSqWIl
FOsmjHxXqUt+KZp4zjQlnsia7bz6IJfKrbCE0e0lehpmw9mbJtk3cDYTBO/tVo2z
JCYu8PFLuQeLr47+RUswVWUj2YHvhVvojTlIMEDwLs3XuZ0PeL0VkIlOH3+SlkFM
24xrcbV7gCJuZM4wXyKy0LayLc837KWJYxk1bWqZh3mnkaWr3vLwAEXRkNXpAI0k
DnanVcg1AH9iecXbeGsEO1pd1pz8E8/ab5o7qwB5WbdZXUWpFASIhT+kTA5/aZQZ
Krm6fB+OXEX3cNmgBuLf81nMkMJVqDW6cjjQ7PJRAmJk4z0Vnk+b+Gz9LEZJbFXP
aLecDy+qCAam1Em6nxcvh07GjMp2pCMEPGVsoXnY7hPjxJalwCFcs04DPOick8ia
zVtZ0308NtzTuHhMKsov8pNjxONatCk0OOz/mclOHCGRW5bsoIpUgkWv91WM07qx
cyWUa32wOx+qEj+qEoJNUuqRyISxzovOVogGGBJtYMT8GWKthg3QKGJY4qC4i0lu
uUb1luJvdrnw1GaGoaChS6+03/3GDwEKN0WGP/UKti8LibLViV12kNe+IJHvTJQ4
fhLyG5i73WNnPOl5TmJvHS42TGNSB8lnXxuXTtZVw6z6J35i+kg2R+KoMBWkzDBN
NE7whKPKKtNmK2pOzY1Ot4p8czVPqePeAFjokbRD/VkQioNLtHjKippdbAMO+g+M
gd0bfYm3St3gtenkr/Ccyq/cIgTf0FC8SjekE52pAeLTM/yLIJ5WKNq9kva4hr2R
eYDUz2Mg/GwSX1lHdaScBzUMXckf3vH7Y1sWwMbUHeuQLxLWcIrv3MBEey0hcISo
ERtWfHX6y+UZN7HIxgRv36i17ra1MCrHPNF8aRzzwuez5Nfx8xCCwS/58wR1M3aa
bUNiuO+SRFVsCJhKb+MMNHZyBaEb3T+XXFLSR6faW9Sm2m1yoss6rt7K2gcuqleN
pe5zbXbIXz5QpxZKvJ2hXvMQiGn4ItAtgXi929s0T+T7uR4128aEagJw2zKSG9Kd
BVwXSRMwebNLAEcNrpRzPbSuocu8VgtgC8+EQpIzUI6JRuWZFZOgiZ7/6qk/STAY
8UE6fYMpWzEU91YaK+AtGBx4LcXoMGd7lNK8RR+ieb+dGvUwCe2JpZ3ywPYhwF5Z
b0bwoxtRQ1GgKlVkLX8SjX8eAQS7xQIrL1S407kBxobDQTpnsLpbzw8Wo8G6+/Qu
WI/G6oyygz87LGYZ43/6g6j+EM1ew55uhugY/w/n4GLgZdFZzg2gI6JZ5v58D4IF
Z+w6T3M+CyNA7imGfraxmADCFsE3nDhbZbvOvXI4X+vpnDgwfkX68NqIu/Pt6Zvo
aNS6DOxrE/oYFeSS/KpjVS3ZG9BzgROZjb232l1CIYAPOtc59KJGYIwczmx+sqFh
N34LHcWttLJeWtEMbwxxULr5tVW3ET7efO6txV91AYgj+tbFUrOsSBNx5btaXO+H
7r23d8g9Xhe9nDFLMR4nGhr2KGG/bMlgX8wm8HFV0qdaiSThnLUBYOSyonEiHbHj
+lbZloM72fJwk88IBZUJ7RMJBsGk5OlzuyAkCPM5XsnMyZCnKVVIBxAkl4VZ1gXS
sEEPq7QszWnoZlWN44VwyS9YQhd550TXaHBHFPnEF+fHvIVV/0aw3s/CMJQhLpaO
5gTevdhpywhcZSyk5MEN6sIJMFBsKPpe+jeZV8D79HtusQu/q5srDCGgA7oT9pEy
vk4QJGpFYGTqKrdfPLg0XwVkBSYb0p10mrSpEfFz6JaDjqXkfEP6y1OKfVhmd0in
V9Not1KGH7/KzW8MTZwesA6a2Gn17p4N/tTdZkLD8aZXiX2WHEwHH5PvoKscM7z2
d1ofHXk1JXNrqP9ckf5Yye7iy9zeCbFyIvbhT1Jsi+e2y38ZvY3y2pztRXQNoHCz
RpTaUXWUDoADgWKHoLCNQAckT6P0jnkr8HB7ZwhCRvTzAryZGPrtYW3+wtMfgzVy
gCoPTNaOi0J2EGfeM5NVygEMX5Rfrzjda1ZrGB2QYiq9wXig3ObE76obt4uHtmL6
Nx42cvUq7ueSn3ii+AL5Plz7dmf3C5s/fYucKaYoz416WHh6UD5mIpW/7EEfHW6O
jFhm6HUdOV68VSwuCy+61zxxqGdZCcgl4HYRX6ANp8jURxLSbKl1+M2ASGaJHZZS
YbJGgJwPjZiLMK0N09fnlzyxlT1/EYUU8QU+YSlV3YLh6YIxGDYczDk3l9GAIQnS
2UKQpPqd4G5hUHXlYWVkpRSUBZw8fkvuuW3f/a5WLGrmwaCd764GgUQhQUOJ9fKL
RJutZIhYrmV2pGz8TDLK2iim+vu2FpICg0FiDlyKAcib9+wd41UfpkuQNM7VoFUA
D5ytN2GpAZtmPNRzaGrbj+MV1fVKp2wHkoKq4NKKyulF3RtzUTJhGGs+Nvw15+7X
WJPdi3H4PhNvq/i6Y2G9KZhDD9I2SvpacstBTvtJfKx6Jz/krXX8L5OLXw/b0dLl
H1Z5oAn5C3zxiczcnX9XD5TT8eQogAKNAld2CuqdQu7xe6IqdlN0JR6FwNctBGvd
m52T9M6XPb+R/FdhhwK427OU/GYCnqyp/md3ccpFPywTMIdOcZLBNAgK28Zngowu
3aMDFh18w22UZyKYFe1r0VOBB3V+jBXv3QbQyU8SNlQ9Wokw/XwiYmvOonpNkVBg
g4ewEWzReBA++ULTkGzYzEj63/ZvO0x/bFLNBJyqWIpgdiklQYPkXyWRGIdUNzzX
1BH7zeqVMYhgmCR19/OOTJrtO82v/SsESBX3cFu5DtE+pZUafpp8r12khva4DlDn
0cRoeGE0kp24aQvIAolcpsDsqSx9WtMRlLvS+yx3ovHdEkbT+HhmB5IKr49g9Hid
HuGG9dYsHReWQ2OVpSOyCpZEOa6B6AZcshFUhnYGIFtXmmv5ZhpuUKjNLudn7CtN
PBABr0VD1MObQvQ29plOsiWBaG76d/rQeFwI+UFDJFc7PWrj18WLQpfXsiBL49gA
1HvOHWZYuu7Wx38liukRpk5hgLLHe87I+a4v/PBlIzCbjx7Z6CCfVrM7xJGHv5i9
r8sOTmsecL+HJ8Gx39oGId31EHP4E1ylcPIILJirzLBos7BuyNAgnV8HfJc7tuHb
p/RJh0R+ougKVkerIRSxk38RFoz45NQCbVcuKSDTNNY3P67selDtPwW2ZL9n4CIy
1CHczVwMmFV3sUWnOgryziDgp/Q6xIIqZ+ZlADHr/Qy9UpEOlGNJD7HPjXFnTToY
u7BevPnOC6r2+VkpEVi/OTKbp4IqNgCBP5Xzd3+9dF727KyslLMxF57pPe5Po8Uk
eZ5Y436VGmFYHz2XBS+EJznoJdDMxYMiYzFj6K8uXOAVYvZaZhnY2XlJxHECpOB5
bL+ezXRgkqYZRJ3uMtNkDFA4hDpNxdS0YNfotcKtvcbBbMLmhO0KdLDqDhK8qANL
JkqsYFw0MiRBgrPKpnHwt7Kp27UiNcZy23wyDMuCmLzlv8//scRpx+KNCYnpnXVc
QsCA/C8vl1Hz8P3RMhj2SNCCBTXEADhINs+3LDxYy62ZTtCkQGT7lDFUxN3g41Ni
HWOd749uLXnxMoyveG9Ej88kW1VU3IGF+fHFrROg2CwkKOICfWa7A3GM1CFyPHKi
o/rmtHjgoH1jjcVU52WsjkVC7wMKZWeAxMearMesrM6mkVGom4LCWBsro27QJtbf
TqpTf168XNF5+ek9JbP+TqD7ILEC7IZKrcAEuVLTfP1uVP2dcS88JOwaHHouvv+J
03xn4klISA8dV3YBYUWDlsJNni1ikbKT0+Ab1Zh7JRY22hy+Eid6IBazn/WduQmR
KWiEdFSsU1emATBcJusP38wgiaYzPO7O2pp7RpnMc6jZvJ8kQvLAT4KuNvM7U5HG
d3kwl2ClI0CLl7he9z9N5hPtQ5Inmbx0bbw1W96jxfEsghhQ8YczFSUTAMtJGzHa
xJBZfIxzwft3iZw93+mum8vE4EHtANzY4L47+Bh4E6O3F8S6+TYs3M2dlDnZJSIB
WMFUakcpHFX3hA2ZVuOJNcuQ0gvcAJv7zDD3VG+TB9aCY57nmMsXO3qyyvvsj6Ls
99ccL+Rt3OI+Sxf5Rty7w1lKQ1NwZrhmMum5P+UoFsdBXGEbCYsB6Tvs+dpEhBbx
FRlRBSy85rAN5A2OxcqiKTpAuHNu7M1v0VwMG1gnDfDnjFBf3tlaVcZlTOKBI/F6
3eiKqt1vp3YGijJ8A189llgfA/43vgp2LddR0gt09qIKUfVkM16c1+ZiONUb4SUQ
pa299X3PnEqh3IxP4j6QN/gvJDB7U9CacdUDWom2++6RSXY6j/ejAH7u6OqqPhTQ
KyoD1TsPl9K8Hsk7B7SSPA0nVsXrMYwdkFCnqxXGw4eS7z5eKH9R8kWAN4UGPnuL
SsjfHJ4c4Avq9jG7DEeWLMlYs7Zc2K3ijDYXH2bzokknbJy4omo1XaZbVt3j3wX5
fW8DJHMD5OBGv9Vlr8NDnsiO2KvMyPQ9mLqQuyxKXHyTsQS/HilKssnPBXVpK0jY
D5czOC7ryf/qnqpoBHFMzRf8KTmfkgJaHinq6Dbi/zZUI8+q3Z+hNS+qm/sRv5eR
do//rzmjxfPZ0P6xQIkLV4ZsZk/IbhqEHfIiH8r6OpFxEplrlswQiXG/ly6hOJaa
OYej0W80YQ6UXbT9TIV4tGwVZU3sQuBpokXRojVHZmMLjzl4bxCbI3O5eqQarTh0
SRIzBOPj/sQNjyKLBKzFyFxERp0OBw0UbPdSYIGbwTBmkX+9JIEWA8N0bVKzLozC
VnVmNi6SLy2EX+cNBuCfpMqG2U2wa1wP7VngBn7H5sEn48T+nSogS1bF+bpzD5eq
C/xTtg0W9OCsW19gxialrEYpedNDA2aUMIbiJc0cHxyUKFnTrxnlDsQKvcTEyv5A
qsitePyIOHQyqfqZTYom0PJKbYgRb5x6STOKxcb1IaKnPW8qpPkL7FgyDBeYYZOX
H4FDraDwelfUUzZ/RZf23ylPUwerm1YC40e0bQCji4roZ58HsHS+tYQErgpOXhst
wEx0v4y5ol9yK59MkuEz9+y8vXjI18jtRAx5KLQvA111+R9uK1feFsqCemg1quaf
qU5LxEUJ0drJ71qDmcdifZixGgSyMgZEq/2RMCmyoF8ZfPLAVUQ0URiW+QLxKZh1
6xbDlkR/+/YEYIMsPgOpcLU+AUCKO1iUt0mw4hjfenQt6PRnOWYQVlbcpaoc9pSX
vNlDSkjvWnFUUCVpmmeAs6MMMKswf3YgUuJKdUFPqDYxOitFSUfw56DQkHKt6L3+
Uux1d7xav29F86AoZ5Wh9Jcb57Rn5K5lDiUv4eJeaGsZr6tpBXpGlLb8xUMXrW8e
KWKKb8udVQLAo00DB5lRoOevxAdHVdhEHXnW16hyyDx60XnbyrwjYcye0f49ZsCA
DNo9ZNO5zCxYbX9ppHspKvWw0gTUFqDoQ5GgT5jDabVvPeTo2urNM9aEd0ROz75t
exp/KdOn4nmHeMT35pPNnE5XaWHWsAkjE6yfX9Yth8oAAGPimj+kRhb6xhZ8JdgU
cqc7muSceoa3cmB1T5MoqVttbgNsPeYfI0G/ID6Ceo1x9XC1k3qbMwwVPDurDsx3
t/YoIAJ9igrmc8tKqwqAUG4U3lNVfcCFiihq2ngjnTMUqOm5xQEhAh4/JdhYiInU
eFe4MIKha8ZWj+zg7EjR5GqIS2gnzESJdeb9907Z61obj7duumI+8oCBAyA04gEa
It5vHjcrMoFFLPI2SGxO0VXomhTN6man5A4ZAcQzTUTDYEyYoi+teW/8cxyo8YQZ
aWtcla1D+zHUTMPCLvBVQmdXYH9OkPWe0GvW0Nm+gMn1qwoveOKLucreUxAsiiJg
i39uOdB5SS1x+bO3oidrysiVhVWGMPgVtjfzWO6jr93AlUQGl1YKnYP7PXd1Wuk2
xzxzSKfw/Q2fwtc4O8FXlRyADm6xK6WgBiiv9SC2nC1LKjRIyJU90vcnSzqUkp5G
MqDnHHgrfmCeELHuLaDQhyNILERjOFfqGSrVsYN4xjTmnNq4dSCkw737zrg7S6qv
WPanl7VivSzisj0Twsjx7Kp5aZLov4dF1XxggY8Cv/N1vzP06AkSw9v/LUxViQ34
Umt42YFgqvbotoum9DWhEvv5BrfSPvny//u5/WKUpbaAoCyn1KNthbCGnoAdxhE6
2h3xvG1UhrRMlWA3vKWnrVS60fYDbp8LfewgAkcE8btzPzT5BWuMaL7Yik6EyQ6p
ICU0p+NK+TUapWxQ8MBBUqzpzKXNsjIXPCc5/lkCUWk9YWdVI/3aziU84NcVVSr1
zv8DdCD7T2cemeP17CdBYKtMsyM6EaUuAHcYTh5NyA+CPMuhWGMCBUIwYH0fl+j2
WSgXBQz52HJjdnLQEeEMc7ONG0qnP41Cnz/7zDMYa6v8sPbPOybfyIFhfH5FdWA1
Hady04GbQEFYbb5YZF0XvSKDmCPTZa2AyTiqH43NQkqOGua5zK3acFt4B7W1cKgv
AoVUxTC1DuTpGiZk5pXcMz2qEmz2UOc4lE37vPdZbWN76TbRC2zKJVYUxYwtUAd4
FXYpMqaVkmm2FjnQsDdvyQmQSOorvo1p+J9hhKSa81Pxh8cGciDZ1r2vdvzNKY4K
1PYP8s+3fWv/qeWpRtysiMGYlojM1s4NdxIu7T3BJ1k9kE9FD1wo9T2woeISmfZ8
eIYIPJpq5UxBAdafESK/nhKOy4Clgf757f//pSnUvb4UjLMh6RuUhRU1A4+bFJGe
Zk2YMq+FCQM1nSagzqtYmFNmzlgC289kTGUCgip1CTz6IjZaPLqUDc/ay2KS9rrs
CQJlwEAX41+lknWh/8JCOW1GgLYmyQ22DqSUz0fIAS2PWnGu5gCqkuJVRfGH/cN4
lY1nEjPiccOyhRqZ6+kIAPo3rSdIN7ppevYHh1rTspQbmJVoTAs0O2RH8wgmdnQl
/5jAQGQOAiA30Q9Z4FX0/j8O+/4QbmshoaIj5avO3EbInu6qLO9P5GO3olNcZMqD
jyZgUoMnZOt/4TWpLKva4aLVS3xA92dduA5dBIl2rhikbdTjr8KhU8B4YQ9mnydn
dgfEfV87Mu3age4/VPNjhYo7JMUdkXYr5KgZ+DCO0GuyuUg4yT4112mYU4g/D3/m
PjmlFnuN0SY58SzyV/BnbueLfilEPNXLQIZC11ceGVuAQzEI+kSdzGvrIeZ+XMof
qRGwGMR68xlYdbfptG980R6ZYUf2k6+hPxOwbjlfYXvn9zTtJOIlYdf4CiT+bKYj
7KJiVcJdDlg0ffWcHYkBiPSgat2YE3qPpwhT7fnKUskaBl9FXVU7Q3F327g5BNEh
sC8CZscFVLFiCJj+ZU2te4Wk3PqUBfuji/9H6GH9sBIi5zVBL7LCSDqm8PZijjtb
H36CF4zCcY6yapBKMiI+PbtUmdl57BuuznwRQIV72A7k+E3eKv6ue+rE8LfsvGS8
oAWWTdglWv5zfhyhsH6AUVgkmOusp+PDedCC3ojwivL4ZrRT8RP1gcvW35AtMJN1
4RO6MhC7C9TI4KbdMR1EcjvU32TNIK8TjgKU6azJpl//63dbyuKdRktTbz2EuY8W
xOW/iJXvaRVuoH5Wlcmcuqw1015Z9NRR+upd3qPxiOBqZrwt6pkq3fh0Xj9SMPCt
8UHvFqJ12dkBERIX9XfnzuLGt44mwnoOggkmqX8H4Es5iEsZLXf9GYcZ6dgeZcvH
O8tCde79NBtsinGgy++8UKUn7BkxegQGE9L1SFZugCexNLd4DDDPm/uOkpko0YMW
x9jaJD0SOWBFxB6WSb0OsNKcm6fqaPKUV618h41ftHxJ4yW1L6PaETuLOdp3j7Nr
SQxHX2iYtFL9Gk01iFXc90Bma2L+2o6p1hJk/vChuSIwSQaNUVF/R1VATMi9ZjND
db2bDxeV3y/TIPMiSclyYwOM0ylQFjd78T3ousFUR1Uo363iB2ZkEAxXJxtOG/Ib
3TSIxtRcefdqwBXTmEE+q8Otu/+crJ/dDKKC359lcA3Vday6YYFpUPcvA3PsqmL6
ai49SUunPjLovuYBWh5MnXfRF5sDjHP3cwp1r/g8tMw3pbz+5dsTRi5gpMv4ZyVt
DC9Q0+BSPEVyUhHqQnLpjxInFJbzgAeoZQkEFpZK8wIfdU9JGSSu/ynprNC0Ehle
+TcawhBLrH/BCfa1LSkwWuOnzSC9TetPajsPCIOtR9f+xwKoaqYJ6nZzH3w2JQwU
7UYEd2WiWZwYtGjoVQ1mngd2JisHq7nIGw130XcWO0ue1J5h+/Q2wws+9lSWnyiZ
fxSdVTmmcZfG4Yv8B/Zs08cYGoyIJyUqN/Vc9jWhL/Pi0xjkye87ZXVKLUMnD3MV
EMP/tmOWJ641zCEDeNROcV7UR/FHZjm4sDWd04RaUc/8h7UGdxdzeVscEidcedbW
zoWLSqbVS8Igpesc2UfPq4QQiJGvBv3AIMqv625XnreK6WdmovXkw/ZOuxl5dmK5
+A4VPkZC5Fcwhd+DbZ7nxHcD5WkY4LlTciiBtaeN2FDTUnMNbR3Ta1AL/KBlf1KZ
/W08ZL+MCNPTgMQhA0tBRkHq3/5aiXkEnI57HS6ws7fyN6NaCpJl4aA26qO0zNy8
9r6eE/PwSpUDhlvVruahvRhOPQvUxyodKZiTPtb1/qpkyeTxeidy+Cuk2FabHimQ
kfrOpvmBE5trmVuIoOvC8zbDoPBi9xo52+2K/WVdEyMtwhnZDpaRrJXcxx8PIyw+
EZamxrsreuvIS3ETLvHnRN8yMzyPGL1BBzUCfHjf6E2h4HwjnjuOZAPkX03TotUv
UVsGLseSuKsA0KsrXzAP9cYWSaCqaSOdUc8Jjc8i5gHkLc/yaYPFUHiNdcdrrAPN
B6Ww4tHq61wMZ6jE8pcZENhAHpjSWF/oJdSmCbZhzOC/GK6mXHvqW3EcnyBZ0jil
l5ta3grjoaPnIs3R72fyvQXIOazbDLn4PlHqCnhA+ONvH3DVQljCHnvpw/Rb6huf
4uLLo8lN/KMNFHF9Umn79qz8IHHm0n5OGf6PMLOvFNA4DVkAPHNWUqhAC3RXIfpf
inooJY2BUKWYSIqmgZoTU5OAGdQQOcKH0dtZ0P0ykBCs4O/MAdqHrQUvtbPaOFk0
vLMBYVV//dxqe7ASFfA4kQt+qA2XKJx3sEvgpSJdmYD41ywHYBuiSjlF5eFUMxLp
YTaRagsTRGxlPnmRPhsqdxovbwt4p9jXX6qhB7+Brzv2V8jtzK7rDQ1Kd+AnE595
CFGVNohFrh6tLJ+PIUjVZgEAi3oJ+GV6/M51IScQQR9jmEQJ/eFR1H1/wSbR6Xf/
ysnzgDBh5+XDSVCETVTQe2hkR4EGU4DMDKlm9HiLaIgW80z1bMeGtwYU0bGBMDan
ZDjFWe+PHCmYCdLcU7s052VAki1JEnJ2Qw1V96pbGv6ZpV+4L1t+mQDvETqRWjO1
jL2Va/Rb2X3wbgbb7LXUBVrnV/VcTC30XCFobRhaL7wgNhTVQ7+3xnsKvO+v1UX1
Y2RbvQABDcUxXJrWCa1EIOjhEuLbgk4+K/Cq5asuNxdv4lPrfZaXXiB33pWufrAg
HBLaoxDFwrNw9iGPI3GCP5kgRi5Z/1KpnoLQXyXpG4cnsG4GclTbeG7GV2ck/rnx
qJllVq3hUUetEgEeqx1qdygGUCMKdZ93SV5un5RDE44aSvLGKpuE1ENyfyBVbrz9
41N4z/LrpAubvKsPRQAwyEUC8jQovuWkVHGFe1tikkIFd4aCBC1MBU3rtfs1HPk5
iVfgpcTorRkDamo4IzMOtm+aAHgQ47cmUU6bXTU3TpQwmsIccuvd8JXELZnemOUM
ZIZAcdeknax3dcUlJeZnRqVY3K2modKJSdDdU2qMo5XV9vw857zLqwBqTaVLdH0u
TmrOCOD3LpnM/98TkGWuVmKf8uZr81mmkBp0rXdibYtoDmhR5+7YP4NFyw/ZdwRz
AqW4R4DLE5dhYB0kQpQTY5FQnE40alD2qakYzLeR9TwSoU81l4iNzf1ORxlC/0xP
xjWCGjfFKHu0DJRIBynmJ/JdkVDMlYobLTX5TCPfdnoNpJ55b1CkuoyfnAqo7jkT
CqSaPxFQcTCN3mQAg20BUrP2yrPJproyOnNJaKhYGSLl1gwu9f1+LozAwESfHn6+
vMJZTeknf1QTLtlmZgzuvFo+Vj6KMshhDdfvLG4G7HKWANt25RC4pAhb1FljxNxR
x5AgyVIohuvhwH3qLPe/IbX53EToa8xsTlw9UwO+rzDJAazKsDTZkfV6M9EejXAb
hzwpTTbq4UYRLNIO5oJ/CmuvxiSE59ukkQ7IV65e92E6qUCNUAFZQ4i5gjplHjFS
rYfC0S67d3HAvCxnQYY9e3cD7uwYDUKC9xXnMZFgE1j5iYoL65ywHpg2ru2DEel6
XgZln3/yW+nfSB7dVBttUlLW/PAcpQYy/iI6qlWIdiIpumFYxZhezK2JDllA/Je9
g9NjT+YHMchLSvGrc4mEV9TRJ+vU5mWdRoHBG5lxeS9sXsqrluasLxMPE415Ih/4
5FgKr8M0vxwKIY4nY1KCQeBKCXm4sk/V9fZ1Ztk+t3590u1w+MW5thYeX11RDhC6
gmLXtnaKdfICuEzJePjBpHKI1tJKFYe6eKGzgAOk4zCWc2pEQWbdMjgpxtX+TCQf
BCWcNdEYNWy8i2Uo9pWfRNkKFKassttHQ6KXSoqzZIdWWni51AXXISz7jK/pa/YG
05NSDrG5+vbrxz2qnhFDGrJQvSOBKtd5YTIYB96WDuiDtzCnnbLvPR5De1FnZ81v
L391Jn9cp6TKJGXKJhIPHJGSF7GPrnCVklMDPD+QUlatKVUOzUaqj77ff7Lf4Url
HoXy65fJzizBgwedg3yks+WYJl9ZU+3v+XWpnaG0BK51+EnfnlSbWOjGvSMH05zx
Y4gat6W6Kw71uU5Jh1MDVXPImI9JBUiJjI8VDva2yiqzBxqgPEBt+oH3N8HSAewr
ell+BX409vFtOoNmVJJibc/R0tuUApIkANg55za8injPooksuEBNTwQalLAL8BbX
yWCqin0WZ93iqj3VLM7UEe4MTeVyY7PTb4l8SNIaVlJPS3lKxm0FIEgtU4aU85O3
KC06puN+aNTDYYSNovQtQUWBLvQr/hTGn/sJYrjoRPfcAVm0I1e7U+PIViEc7+8Q
v1lvCmHoGB9vLnTd8Rqx7mCo8pfBHCeE1MrhDxkaJhLbOpvdtKVyN/I4ExWK3RcG
UmrJHKfe6dRNHw1SRzFrDw5iQdBZ0NiF+8nZ5GF/iGze7oQDbTNxKSPTZaVXQVxR
VhJnQo1SBILHpaAWvzyLv8VW279w+A1wL1P26bQgzugw7i7bBX8xtfLPIK4erBQ8
svZCAfH9OmNTpvwPIu0vQlCIBiEEFkz1CLN9jV9SEoU0pwtkHyeP9x/CX4Efifqc
+Ci1KZAleA/uimI33CXPHxAX3RyaxhJnipxx8AG8B2gFbRGj79j0RY49CfzyilWb
HzGyFohucVOjjbhoH4HwVDo62dEaYiOxe1Y5q+VtGSYgdjeVFMfljxw12jkEmqqC
XudVrzlJv/UpfJP4wwwe6LlNlLUCNQaECBImzv6DzkbipIDjAtLoXwPFk70phUFC
hItepJoTp1gZCBzg6unw3KA42vj/FK19HNktFuW2OJ5KiNfvDQapK0SMlSmcO8Vx
/7XMHx/2AjupZ1S2ayGbQLTvhdK34L3wUjbhWKHUBZmzAx3PHmRjVdI5UN7uReJ7
DAVLKX2L8oPx76XCwJPGjpxUum8mE89YiUKCug8F1pr+OI/6cW/06WxwnCaOQksB
+IidFEVfT/X4ALcMXFkROwLO1Z7n6kjny+i0ziIx+frH9PFk2NH5LJ7QknWKXGhw
JEOSd/HoLEGH+FsZ7K4kd4Qd0tqlISLfyG8hLIqRJv2lCI9g7chNaCfuYCXr2C/d
ZgkT+5XzlQWRm7Z6YErZu5I0u63v9gxJP5yjeCBtKEyA11nXWtP+LVOGKXF4ePcR
8DPrmHP7eoyD4yWwotwNLU32s8YG9Fd/T5RHt4MxbUbdlx/N+yvwNXNmGvUYCboz
ZsTppp4//80YTiT4Q3L4HcOS+/FscdsDvljexcUaHmjjgXVhfUEJrIOPSEW745JD
R9sUBWKZMe7ga3QjofTHkHqk5TLPh2s6a8CYUU679hrfmXnlOjeSrUAGBrhx2Q6A
/H1XpW+9CJ+lv5e+tZIB7mSDq0EMJTW+aZ46gSAMl37TYwJVeDk/46U/JnhDyQyl
yAfsqbx+R8+9Apkx8gqJKzqLTxhMt1zAy9LrG+7nH/g2Gb55sciJSegKyNErNrJT
6swULaJNWKLUp4eTQRNQ6p0SvLxiIu74Yrw/ML87EZdRgq72BlFVFjce9W/IyYVR
TDyI7whvDtA9o5rtF8bBUIPIuXM+vxI7Mi9ZxeIcU+7TxMORGN050Aqccwvz+hzL
RlOTzJPzcjbEmgdwsskLfmDsdLLvjnXbDj6CZT2q/JxdBNo0mk8dVNhpkn36lEMP
pCLLlMdCmx73iigCGgYQ0zQEDLdvVZX8frVFrhG6+6tij64wI5My490Z1UNeqDQy
b9De6AJmBBJ5I+9ZtqoFQX/NFjC32RMMxeJIQ3eb0jbRZFh7r/dU21Ltx2eO/Lv+
pPfjYPicTE8nsW8nF1FcBpcikQaz6D0g60W09pIf0wwFXY3kf2SidFdJcmeY/kiu
OYED+PkHN0wH1gwDvXF2FVpcz/og6lJRa0T6Wd04Od13/lQbBzwedyqz57S08BUx
4C+2B3pTzT/IUxBZ11IoovHht2cF/czTncOTHs1jk6y+8J5qpyF2JNywH19Iwqzu
8mJ1l7p6tchKsscrnsSv5le52NNxyTzyC5S/xFUYgBMaPIIy5xKDzCakDdz7mohd
qO57HETwsoY4BSDFocHKtYemIxzpknDOmMJI0fsB77Q4yJxlAsn65VB5kNyJdbHt
UFu8o3Mn3bvSc6qaKt64CxyairVh3Su/BDbOAft9iQ2oNCwQ7gxRKmsObvyCXPv2
TUheomgDvrewcNxNe+TJLJTbwa5sv2M59iEDJ5sQec4TrKPKgkyEZ/zqPBf0oZGi
ym6Vrwj2Qushyp6MhKcAUO/tLgNiL5Z0DxlzGMHec/gLw8Yg7Y28EhrFU9ImDBkk
Vmm0Vxy0hWyxqCFrPfc1CbhcmxvyC3tw9JYJdcCklBtQzYEmEQ4OVH186HHKgKak
enncrlo23RpJnl6WXsuA7uOUSJOIauPL4Wk6dReKGol+OIz6Jj5xJZejbC6Uyphk
hBCNTRTswPtMXAeadw8hMa8JqI2tm3Oomh5MUreuRuThVU9uO4Tkh8i7+ZkFCbHN
Zn474czo/gNy3wrvX/FJB10VcPGW377L0RNuHtW4KyFAGH/VY2fy7twTSrigOiIg
3rD6wAQzLk5qX/fU/CeQFmt8/Rn0q+eaajo11njMzOG0gHmONQxV1Tn5PzlQpYRg
2v1rB+/9WdeR+52nGS5xT7ST5jHaGTTZRgEN4g+kusHWZjOQZ3OEEaYWz8O8S29j
XRiiPwOzMawDguyHsbww0iL2KJafz1qZI4AB38xaH2eMl9q08N4SwZ7FTVxwFQco
t1TnqwQbAOS3EfLI47MBAOeyIlMSFYu+qFhYgiBRi43tb/dEav7zeUcvvRR9a654
9rn00z4rsDcCRClgYHiUVNMiycrtX8sGCqnP0aNSqaXLJdGzDa5VnSBrty9cVrBH
Yp4n/AydBW610AadG/xmNRLGdVJXeqir6yErRGPcKSqOP7Q/t7LZzj31dGMAE5mu
v99RzC+Hg7V8sNApZaazDvJIn5w7KGbH3lUA63pgHcnwxKkUXx01iUSHi7lE7t5F
Jtc8BAB9cFPZo3t5qLSRZZQLyOg6RstZJ0vF4aoyrp/UfxbqQZz9O2QOPciLwCGD
uKXstaEng0yxUinRyNn4f9w5PQqbFXVbUGVEtmgUZU79+TI9/cesh/4AG1mxDnUF
gqr5GYLGHqGrdLm7rY0Ga1PPWfoH7OkWXWZ3ZzNeURYbwFlI0yMW4WA3R4F6mrQA
ozmNlntlQnSlgsA4e8r8RrM3iyNaJsn1wA3B2BhsSc4kO89pbOEHTOp1i9U5HV08
fcAO2m4rjQPQbSWtkU7zp001B0jDOJckgizSHmRv7X3d8DxAftP+LncwuInoApZg
KoBiPNiTOsglCBNIMkLc8BDwIQNVBrTDCleTPCqqSkcY/z0SGZI88Oa+Dj8P2iF8
xEwhZ0ZeAaDHiimVrVgdwQNEqzxRZep/CuavbGkdCLMUXXViQWGFDiDeUQhqW5TL
51SVIAd0Gk/B31D6aah5MqRRwZsOXpvPIcchr5tghjr+fyPEhKflEIAaaOZnNUh7
D9ON0NkL+jczdZb6m+MmoHXeDQ9H8M3wQPTYtXnAeNl+EZAyTIdjjmDnfSqynQ/+
aMwL6HI9iTfXKX/3ZTjH+kHUYl/KW9UgDKcwmNzb/jZUhJnxHTn68Bcg5DeqVER+
rfKSMjYzhYWPpn9Aqxe+KzROYsQykDCq5DG/0jkY0d89u8SuluH0FMx7NKwTa5F2
ocHocxyhHfCfq1IVRS5T7pPkUhH+PrQslhbkMndhUBCjWHVOGu1tHnyjbBsQn1++
OCINR+IbHYVKSllzA0oENX4EMvcExC0PDUM3lDhnXPTiYQyrBp8pH6A8MdA358LB
JANCcJUNq3RcPsG7AxhGJ7utSQSGzq1BXI/d+trF4EK6la9vE4PAAMmjqR5LERuY
6YgPAldqPGYNiNvnIa4PaodW/ECxXBY3pc+3lFI59ndmZzN2Rgl6G4yW3F7X59Hg
aXPzSLt9pXraZKaMfOcgwFCqVGzDlYJmcsQjtiCGSajxMCWaS1Jrtjbesogyh2lN
S/rjliXHd9urED/XOPciqk+FgZQBKoaAQcqC8XC0NdsEHA8aVd7d7w2ke1bhNdqH
wHItOyPhIfuNUC9r31CbEc209kVB09KXNR5JQKEKKQPGhEQK2BmmMg5Kid5AtE4v
QPgvzb2FVZTpWUgdby11cdgF2K+vSYUW9EMWX5KhlPA57eK4SmpemwVa50TlO5wl
0IuUqhrMmHfKnDmctVTaCB6m5d9YMLqvSBq08wazNcRBtPrjBaxMwlOwvsTd34Bl
c84H7+vii6k0iUogRsN+JuoUr3sic50Zd0lrbqVMV/NJCwQoaLJ3bf3V8BMGUOli
608+deLSZfHVRl3ty5oddJ7CdWLZOL2IfA7mMsCqfbrB2DxzyNOh6B9JjPAdSNKT
fJsuGolA/zfT7tzkgaiHHcTQf0u+lOoIl8pOgRUF2rI7Dj7QWNAEXLpx11M5hg+r
WShWiMsmFWQsMdTxdquUHpjqVqyTGt8v5BiIN9Y5vskIXbjbhPgnv86+b6vdXWX8
OiSxLh4htoHzzKgzB/ma+l714caEPmvlmi3mWn5+8SATpVw4NxuVuh44fwF5wjYB
1PS1Y5DusHM6IR6Z8Kk8jhYla0q5ulOVTomfO35XZUo/LZmvsqMpkbB5oqTgpRl4
6omfNf3vrk7IT8kvEReWgAD5lQux1GJUr0VUxmvMG/oxo6hmuRd6VDiMcSzIpPe4
9Gh9Ymxz17a9f4+zd8f7UkwzguOcph+2bC19UJP6e480AVoqGDF9nJ8A9uMf94Po
TPZ1dFKJdWcDx9e20sxDfxL3SdXLz3b+UxQKKqrsZ6ExySgtlpUn/7kFr1G78w79
Jj2BizpSfff1kcp0nOrgI1Y8Zo84FMkSj+iVP1REriSz6uHw5EjK1VHdxUDeMnJs
dKA1rr843qHTVNA9R0qCd9/uakgPNq4adVLf+lc14JPOUhS0ITNGMNYEL2P7SES0
olmMIr/DDa2d8G3YGlrLEw8cKp+Ch2SNG7VgrPXDdB6MK/GCNcnaB+1Id2tMXDg6
ECxHJW4rOR0JkQ0cemsmv/3OmCBJ/OcI4ybiVwakz6oDijZqBHhiG3feFqgviB6j
ASmajI37Y/MSPg1xQbyauN57eZFpFJwLS1lsNHufnFZzhyOc+FDqwUOuAMOPxxEP
sWJhjlTTmR27VyLTkFNYzpwBOQmCCBXBj0zQbYglCzZjq9bxLnMTdc4ZlMfnelei
LHUSEy2D8D9wdoKw6vY2RJomqEPmRYI55jBRlomNPl2xrP25V0gX8tdG/VqVdiST
XhTrf2a52fO0KvycqGmfAsJ197upbYlGvFzF6l5lhJ9K9R14XFl+pBiyfdIc9X+B
O93SDykh4XfyVmzJDHYhOWZ6UAH1hPovjmS7Bt9N5W4d4lzeF80HXTndkVfRedFD
MT1P/rc1wG4NGBh3QU3M7mc/u4ysTODq52TFeX7g2/luhkjfRVeghx1Ns6CqUGWY
jIqSgHpr6V0pSj+R7EzAovijwBn5W74bIid+wHvuz9CTeYtsRUCOYTzH5d2jqdVe
ISgnG4DPSdd5EpmzLtRBDdfgPoczZW7IjKjwee6Zji2gQlb9nGAxtyD2K3G2BQIt
hpTCjO0VDcnVol5jU3pJTDKXt31pfkgDFTFUI91ra7TFmokmsvqfK8jbpD+mzzi/
mrUhLC9RQ2LQb+k9cjYGj36wcaZ5loxJQet9ta+krxuoG/NR0q4a4jwp5FO97oLh
ocevOnJvIjBIhkF3DBBSpwCZ8BuT5HhKoSKK/HczSsykKmfLEqu94M7LZJhUYDV8
dHmXz+OyC14xFmNEkGy16BK/Cy7mxMcjZpVDz487em90U3mx31XK/fyW5gopUifJ
t2ckfRD+JzJlHD4babAiYG4KE0HElBSskhl13LvfaJawBKmIGdsxkzQVFghhiNJ5
e1sY7+NumaylA52kGEf8j4FamZgWyFGcSdnnoxR8MNE+CWy5mQ9TDA2+S3e4nVNT
fXlOsXZddx601gzNs3ToTrRy1vrBlOo8Ejosb4mkmrcGlzK1IuXrZwO9LpuFotT7
Brm62G68e5k/S+iq3GqQ7n5z6qNu6FdP/4XMJU2cWZytv/ERpMlYnC9HzuzhLw1f
OJ7KvSP2lsOhCmNpz8TdEhrz2TUyjNqc/8pneZWFxHGOCAvOCKLrtOEPD2QE62tA
OFUAjEI6F38jlYBSmFrEtKZpuUQzZfnr/PIlMT4SzTftNIb+/2K0D+jlxVB/9XtV
onvGoY/G5ROIcfnt4TOdhEcH9LKTv8TDnaiUzBxNgY3iyabl04bj5L7xXG3gHgUz
b/eeaJ2vH+eVjxeWQDSfV8VvbYdBl7WOvv9VPwi/eylhVij/7z+qEb9te6fhmoex
2MvKDAFaJig7C07GpA+wiTj+XsGwKZB8P1hNRUZnIvVHRZC1A66cQMvL2OzD4BFJ
tsoQoI6lXnYWkZGvI/j3Iu0axHmRuEkyv+4pdT3L+bNF4L9HSyYSg++9cSUtI/bM
8pJ8zeIWXvfEmKFRX1ufqXbfuZXBWE+o/yYgIzPvsJqmMJCGTf5OqJdgnc2SQsr/
6dSaxHcFfx52kgQYxSH8FiTjOv/LkT5OedVM2r9Kt/5V9EtAC4ong1CvbZO4DoJu
ypKm22xqGKbzOO4BbFMYjd512AQ45IinBTQMicUOst652lRrP5M4ilGlh8bztUbN
U/AfcBVe0P3dTteAArUB/vz+Zio10b2IYhhJrM2z8T9wdnPaLaVa+h1hSVp9w42X
hrDFEAoIm48Fmfe35DzCS8+5y+C9NQCgGQJhVQ7i/adSiCIHK0hUpqfcL/DHVsQU
xoCNYu0UG4U4C1ZhntxM+cH3aJP7JGZZ2YbpmTgATeYBI7ljYLaOdzDN3OPpU9J3
gyqAB2KdULMBdWFkh3HDI0POTgtMlV4eMq1gtZ47Lg304cG+ANRiVz859b21dN19
0K3dpw/GEZBcgwtWhjm9YuL+rferJah5vaKmpxaCNzUWcDLjRIYMbgUNWzNQWsNi
SJ9qN6GmKtgn3VUsaYtZ91y3roaqJ7OmzE808ZgQcU39K+NrjxfYZm85PqviuNjD
Lp7fkbXTOHpgKzmAq9yNQLDGxTLu82JuaPZ1pm8GOHf12Fka5i/kT5bsM5epHnmt
jRmSzjvnQuokof1v9uFrvqpp6YO1fUJfDk2hZeTXH+3TrdIl3pwaR0gwAtGStUFX
AIA/dM75njF5udYsufT2qVHACfOjnycp/MwtxkmnC7bEhOgBPp83UYHm6jsJewtE
IPYsqhvaQt5TNE/Jsy0cSaD/0WNatjeM/oSqjK4goO17ebhS1U/uPsQgIYV+FQFf
DNWxn78/MNr0WYa/WzCW9FZkkCID7+w/7LjFwy6HOV/A26/NzRS+OHxibA/01d4a
NcTM9iDpgAnPgJ2dBS3ty6LBTN231fkAFJmf9OW/IQQz8zRiGvPoqkU0Iy7IIJwl
x0C8jd895GyR1KzaOUM3kVgTaHO+sncbabFG+pfSU3A2SC48fczEuhzWvSNk5xKI
js3AcZt8roqsL3Z2fuXOHwVACDzAOb/e8FBPYKI7WmI+DvOfK2kz4whSaOEGtQgh
8FJcz/0B8dnnJPPfiIJtVtpRlk6ojcyHssEF7s8iXAT1SQE9knKAXAlE/wwKyQN3
vRZJ/uJxOl+90+OJq3O9DbXo7blGO0QPtiXMQGTAJ8Q++Jl4ATx+gOtgjvAXIrOG
q0ZJgtmUkUhCw8sS/2tOGXbtIe2MlcZ+Wz035ZIM6ZfmIAwtbJtaTK/NaDTCIyR0
yvdaRf0aHgi2dDBYhA8I9i7Z6tFPCl3u/4xcUIkAvVmmVN16K/rA1LCA+YmnPyTV
yyJlXj61SHk17l/y8ynLrqp7sbgwbXEzLviD5Ooix0A9DWb7Zwv1akpfNA8Kbkrk
U62rjEjElQzzrBo00ragWNgRO6PoBKLTCKjvp/8QzwhkfTZ9Rg4NsKe4LakX53EB
C7aOQaOTlXPH2VOZOz0lM+cZpFV7GYE24hfSO/xLkTl7si2LPEzVz9I53fKV2Trt
uDV0vz0e0s6pXpmqmzLAavGRvWgBPRLavsvbHQHr/2/3S66bSFnxj3iQeRXipl/v
2WCQxfhpFhvy0EmlkqgFnq+Q3SAIlz1bjAHVE/PHX46MCZG+MBz6W1bBAsuxrWwT
iVbT/kFbk3clFe8iSU/wnhn6Y/8nDnUMQB93FDOtDlBe77Wp3Kr3LRf/Dn4gAUpq
bn7Pzdxx2m1dQjxSU9K7fKvYuRXCKsiAbILQ5QTx7aYeBjHNPHcY+HOcNiiv2D9Q
j3n8CEmxk1y8QZOsoIWNzGmDiMMjLZRYHlbcLVOtt1mHG2/ZvcdqxYh/LfvxETS3
ZkdqKAuoO9Xl5R3VAdEVJ2hvmQxPGTkZKARA+G9mUSD321xL1Gw3kglaz9S8nl6b
9ulUaeMV3bm4gqyyCoywn/H8OrEVlQlxE9j5uMHLXDlxPZScLm/gnAIvAFjHVBFK
JhLMxql1Hpo9AykP0mQazIW13cgezZ7qE6YggXBmLCXdJcjMH/hXLclM/ppulTKZ
SYx4SSUQbkVOsEevvafsQzdRuFK72itJ2vtVJs+r4U9G2yio11+O+kPyUSqR7Xti
RNuruxxl5bfEjM2OAuXNQ/JDfKJ0HaJbvLyX2aPI4fDmNo+a9g15ExNwMtU15MF2
j8SZg6FkMcoji2PMoykxPsA6jfdabi0vgwXvToaLGt7QtD3JI6xDcNmG94Lz0Ypw
ezqSdnw9DkftH6XtD/LUxM3s0V28ZfcrpY1OW5RAEmSyMNX417EuCJBDmgVaXWkx
Wmpq4GIqybOtfNQztqFIpfiricUr+X1+W40+due5OlVxF3peD1otQqSucQtqHnSG
t4w6rqhl+1kCub/OzmP3d5UqVbgrKhKQOIfco5R5UycVAVpAbSl7VesJNZbFukdH
tFTpt1F2TKhTILxUHQtKCVxkY5am/KTWMEd/Oma6tXNr3lNtjXR8iFyUnmGehrhv
JZLOIvNky+qkgXNW0sRnnUXfRzCjbGbe6sSNmfk3JGhNBlnvoRxAq0iyKgymHKVq
q0+8/+ly6hICo1g3b5fW7nYwgXkNspAPWIR2jYJY4XE1NAKzwZMy/Y/xLduVDsKq
v9jez3ZcxeLA3ovNfd3brDSzUwe/43cJNGKyCcWwZdYcCOkgyL9CkETpG+6iVdy+
iOcyhE28uA3DwrSMbXBCv+vQDDea6ys7eNWAVsi32r+7nvhTCAi4ePzkxiCIW8ag
lJ2YE+sdUX8rkjy43jHSTIsdIsXMkb0XfD2jGkPU25CYXz9YhvZUOCxxHHDCyl7R
/vXLktGSNVpR6Qpy/IHoA4Swix7tGI2EiRZMIA/1ELzlsji8rtee1PKHrvvxCPoM
mA6yjXJLJYuqlxFgolzqu/wNekZzn0MPSqQfOBv8x6DxiC9oRZ8NbUt+OQtUZwEQ
JZWefPsSP8S/M8b4oouyCAgpVyP3C6F6+DD6zO+25QgpfdFUpswvDAT1ez6GE0bn
I2Mwwqt3HLJSbZ4iQseNAgfL4Vk1xf3656G/hdNcDl1uvqJKlz3ZMakY3tO9R6g+
FOXKH3bpSjuGvSgMzA4HyHpi9Oa+v2HnuXtkKNHr/Dx+6jhRJS6dsLfHlpK0v5K+
Z409poJ+W0YMZoZ7m52tkzq/ke9aRjtwSFQ9gKTv/deIesl4wiyQMoqq4YE7xTyX
quFWS0sHZ7qDo3ceOCEkrr1pnXgQcIvmFf6xrrY72xEZDM3cVGIaFn+B/4q6F4AE
7HNwUBECZRuz/jkL31ZTP92ArTGTYNMYLL6FoXVthOJQxo4GKtFaBLpAOVNWRNVV
/AsUOIkdH1+M4yiL1CNUydOgfxbpAEuzKPxau7An9X0qlfobpHdVDWPhdZl4rQcJ
vbLmGmCF+WoABY+uhp+3ehjn2FrsHq8qD4v9nKZck7ein3BiunqtQoTMEpabuBRR
ZGmVLKeKbCla4ATcvfwnp01lLM0MRkVhZta6YDBaojs1R2iDyVqThY2cga2OrMTR
hiKM2wdpFiDEcOiTOr1T4nNYgmUY6Uwus8YUEdGaTlU1tGhP6anoLxW1cqV6TULi
PJJjpnkxK6ongkuOLZNVoh8c++zaHvKTtrJKgv+9LTaqiuh5s31VI5UvjiQERZ2x
1TjKpf9oK+VN69ZUTPppaRIFOCgyTq/zpTOoFdJ842jWquOcf/ajeAvV1ph0WaiI
IDwQr+Nt4qcrM/q18axwTkyOvAq66EI7TNcwn+V+2114SyVSl95Fh1oiA3QLWutt
/DD2stV0hYF/cd8imEXf7XHzfwnUCJhNUnq7WwDivAbr4IsVO76tLAeeheEp7tA/
OL5wKuWAa/Gr6oZFGyS5LvyAPTH7E7VUBn2TIhg5yhF4EDILiFnw3A351Q1YfCwt
+rMU/+QC+KlRi5WaK0ww627brLLmjw82nRdjPyKBdlLBEYfVMUkQA37rri3bs2IV
Moclcq3zdnyM6xH+w/0V01P5Ne8hBV6rQp1EonHKaqOA56xHYWnyn2KzqlZeYmIC
noSXCL+utB7wENcPJgbG6EkP5IKXVBljTWKKgKIAXRsXGOs0h1Wj/kij4UQWzYwj
spklKQ5QbGAhZg/42ObjhjIx9J2bse+klvedslpkxZbjqUDBPqDq2VbeVcSmHxUj
UIKe3uEZNwf9XKxe8gy1WqHCeboBDdD+HjKmB9UCJsOP43gq1j6S4lo90k22hOa0
DHfT3AypRRYhC3mNAV+Bzg22kWQuAX+DwOcPqgUbq21aG8CpiwfL4y5pz7HCMK8S
eUyn9Lk7dCyaEGx8yLyKXg3HD2ABrb8tlgLXxRRNxv4WS19ePh2Kf7m8Jlovrt64
iVB5C7S9eHtBtqVk4JVsGs0MVB200v/k/KZ6Y996xXNWz8vFORF1O1ucM7ZSsqeO
Y8/UhwGQdegLCnAp8tl1tURb/7vBpT4blzXq4fFgI3LLO3A4Ws4Zwi6RkQKjb6w8
WgfujCWEDPU8RFX7FPDMMaEhI504w0qtpMdiMAxafFbJWxr1YTwYafGMIBpSmBwL
qGgSyR1tyuAjZBDUzDUah3vnwhVsT8ROedwPqtlO2UbVFicmi6q8Fhm4178H5M/m
tKOmqtTzYlbKqPX1Q7EcS2PNelFB+sLtyf6UKnf2tT+FqhHCyZsAWCSmQtbji8sn
+2i3zCLTnV+C99OcqMCUd6c5sSwXn8WDUopDXXvw4uK2iorjCJfdNSX4xp5s2FRE
kAwOtPfZA1mE/UplV8OVzNuhlF3ae+yxggUrb+7njam/0vfyqSTQddOtEChyO+fW
2MyKs2ITm9ij28XeliH6KfcNhLML6Xjl2Anv/KRg9eVCyb3AnCBwt+VhKHbSMWkC
i2/wPIDCrwAkGz/XUjTIo2TFzVgcmVyAXtMkCWRqaCabD9tZiECxe/ie1DBSMDfd
eUs/BeNrS9MGvh56SJM0d/ha6hZmqybwR9OHoXtEbUHR5Z22+QZAWhSW+120Ao/B
gSWTmUp7kGoKkodXtPdnsZ2YahvGFA4cVCgvTnKrQ/XlVTSQeQtGrc9sGp8ksul+
pxNQG+0HP2jq4Kwzl1wIcshCmIeVRrhDnM6g5Cmx+RuQgfXbFPkYcW8p9KqvEFPX
alnxMybAisUdDFNkVNFjrVAhYmUy82YhMrJ/BnEJ34XCRXPjCcZnxix+jg1RH72x
QPEkLN3NiZKGDG4wXiTFv9gVpi94GaZR4I4QxHLSkPNb0SZy4elt8gdKsdS1yfjN
MNfjQMvw2VoRCm2vTd8m37RxhUTwGMze2NjW8doNqGoD8jpAQ/qsrL4XJqzlNBU9
0OYYks7PBjORwgQIKoLylqYfLO1eE7sUzUaTo8ExiS4Xn9lviaDNjZg3X2IABs5O
RgS2feM9hJwDauazKk8cMFZJ23+LCtcqxqbKciCIkbQx+UKqyuIlc2V80AVX60uf
t7l2PHrF1ueb+ngaib+R1OBzP9clRprWz2wEwBoSlyeHbBN4LTusMOekKLypQi7d
UXzd5Dd5dXS1ddkN8BATtm5f+VRTihUlscLM77YelNdesYyWmfphlJkoC99H9Fo7
Eqp3pmIbMaQgsMKTrN1NHI9m/tn/Yg4wCn1UrWc0d9hzWx7CTIyC6ZoQ8xML4xvh
TfbuKEKhFqtsbULBHMxoAUmnbzK12ge93jpFBzFSL8g1A4cJ3HvmWLUX/8v9qoZf
m6mmbrWwWqCFgFMItgAfT90OkNBdc+6ewA21pwAM/5g+C3yr3+0T4N3IQFH3rpoF
OANfPQ4HTofjlOLW7rmYZNu2jF2PCVwyo9a0n1mqCw0qY/1U1Ud86pqE7/8kGTau
+4ApMHC5DSPpI1bIG1w/m1LiFXB3deOYSVqPc06s+32sQd3HdGtxRWm/Qh2UqkoS
+4Si68EgAduSebvRebYvVfO2MotGBYeH8c+Q8lgB5R9RMIijAzCBjDmBJDHYkt/s
hLy5MhNhmZaqte/2umNoApyqvlT3lYmD7w0qZp+WmMlp+hMaq+cjYo4Box9eoN1S
GBX7FZN2KxZQOFT9uyK4io67MKtZ1qD0E87XmhonJhzxd3f4l5YoROhouSc8D28P
mawXLN/0y1ZNFmCN6ASNzzeiOwFrkCZjz0SXIPKR7RtiC4Ou6h1E8m21wQPT1ziL
GzeMDMQlaSaZHOd9eGzn7sxzfM0Tju6rA2e3+LlUiicHEv020/FBozG93Yh2DnhU
hu/ae/KS0lqJuQTra9B5LfY7U4yVWYZ+URpjFvop4fel+yMmtgowGNsnb9U0ScJk
xb0eU/BAPn9/2jqE0Nv3eLKjWJvHXRjb9lMk3sogLqGxk1TtGn1b6rDWYy0m7CQS
uCP1q6dpUwzZh0rp8l9WExFvDVy5OUVRdSbKBo9dJTu60QrZxFYhg2hhsBFCtfpl
UtypvOyjL1B1epd9Y0yuR5o5AXQBvNtoswv5TkeSkKhyKU0+xK827ehBr/u21CUl
5Zj///KdjTNNQbGfLmdnhLbwSY/7+WYV9I3PrIoVn/5gOSOkrM+HkOM/uqymzHf4
VPdjbAQ1hEbOX8CiHl6Ju0w+NT9LzOcoXv3hQeLuwEYUrsTHRADoj1+gGcGukl0B
p8D4JVjTpBmkAGacY023x5M8wL1305NsolipZte8okT8Mdx5PENd39Xp8WA6OuK+
g7VSVqQ1nLNGB3owCj/4lpXJjgg4RxwOk5f+7NbCuLBhzaLdaxSQd2yGz5TFXLEM
dodebUwLMnuyicwDWHl9mmNxVyU6yP9ZAoCjgQZhJFXl56fETcQUjSysoMupmy/C
kMsfPJfugskCff5I1Y1nuwWGxYiCARxGi8xnqw4NkTvKnYJcfbKdbQ2G0KDOyjVw
pdU0qVeZeqJgdk7U5YDyoGYcNWjnOG75FzT4CeC/RdU0OKxXvC9xhFO4mOrzT2w0
6f39+ZtS7ySBHGvIF0VIkwukh0Ue/DKNeb8gZZ3ZxgfadJb/7JRmRl6qrsoCXl1U
PcTh+eXydKweAoF0vxTMyEBKgGDAitGpV5Nl6Nj1jJdq6IKFgUYlIEOMYZmv+HF+
2wiTlH6PB38ssFFx356txUbWbw1KWYmEGP8Bsoc+iCdN7G+RGkKMp3nKR/Buiv0X
BeFHAXA0RWsY6iP0k5x4BaHO1dHnDgMY0QxnNB2sqcpSZKa1LPEZoM2axkzydfYc
nMtNp+Nv4453uYABRmWi5zbPxND1CiLBuWW3D5pM+ZZDiR3PeQPv92Z9Sa7Ba4GK
+TQ307ZSzVUZ65aN/HdUw2dzH8R3Pe7vaQYAlGX/2ldocBZl3/kF8EXmBMXbs+7q
SekSf3j477g6tne4wZqUgn3XnBQna5X0tshjnUAR7YQaala1DV1OjIhQIJefYC4c
xP6K68XJ1BWyWgM6APiX4cNnrGsK18DWcedk76Er7Ly5Y0W69NHbf/pCsAUSYzBM
F/rE+9mscm0oUvc0YWuOTJsXlbzImqo8w+cnIg3wkXBaxha520xN/kLYiDu69/JJ
DTJr3JkaMJS4uN2xcP9MAwhhDSWxlvE/L94XmEFA1x2BFDmHmjiiMtixaoDHQ58D
d6cOUnc21h4Hee67vYKGxYxYzj8Lox30R1NF0ZTKPvkO6J4DGsFInmIWzJdNCjmf
zbTAwkpaSd9Zehz4vE4I3KKSRHY8dX/EIgC3NObgTH8jrWFQSapIh84KtwEwpLD6
QlpRxXI+hnsXADeUM5ndLYkXRbF90TlnDfxgZbTtSpmdiZbqlX6oJrjfnPtM22oe
WonLi/iNwyRcZX3eAPnNpMi+771p0ZdsoUjKeI9hEytDmdsm6GLj07Ae4Ik1eaNV
CX1ICQ9Z3CnUreGqnpkxvOK8xJmwzo/Sh8oENOvU3SOiL4DO+mge2UvsyEnUhGDb
sSQ0fRZmi1sHuNu21ExAojup6AbywZ+vURYk6gv6op+MyzYLLj3K90+27EGToEv9
Im9bVk6d/EcFw3jgSiQrtNNY/lj/ROnjPDawxLzJT7PY2PFI1+4StUEo9BwG0rdx
z12MUQh6rd4SJV2WY2JsL5Y+QSs47uLRR9v3vuAMIeiovfTSxhNIV5j80nJ1PXej
fRd1rK6i+iq6zliBwSk9POv8dYs6Y2EMCDKV2gw9yHYKNlZBUmRjyytaoBuV0znD
IrnLbNFjioIsTKKow62nA7BWQAi5nxab2R6/uq3RcW1k/UB4XLj+5eZwWXSk2S8A
LwF+e5/A+nmWdI1ZWiyMCHCdohra+oL8ZQhZkiL+Dg9ZJ6+wPeXuAhx3iuSwbReS
XLvXfhh0IoPMOOYJ1PYCNrjmFwD5VDbu84gHbF7gY+2ZiSqHsn4TT+lKycK3pVuD
gsuHF1kNK0uIdrT5S7/l6meq9la3znWqfrzXA057K+lN+1eGsiQHaZx5TsFoPBYL
dG06TBb0kGUdcX6U+Yga26uLwgInQF4o+so3tbXT1QEj2NiElD1Unrdnl+iVqZsa
RjjiMY2yNwDDZCWrmlU7o75Via2vHpsBK2usBTeCWTC+k95V0ESiaxN/x+c5vk8s
d+uMiy6x4LWsxyQiLJt8J/Wq6PxQNPOmdI4WfS337tlhFb4xugS4zZe36i7sX0Zo
ocFKSzNymJSvuBmwXFjNtSesJDoDiC7RWxvV1PJ9QxZuYdPZOKuxsK/fs8G7QCMG
/2NVbDnRnqM1arTSQraFlx1OqWPuLMb8E/LgQ4qF5UKs5odnpNsNILFwnyNkQtpm
Dl/2lUEbHpOJxKAhAEUPSAAGgCpNQIvmOFLGZ6fcYQyePQTHmk8EvAgxrMk2rVe7
HguZ6Xo9AC4OueeB+uGqzrnCLlimATlp2NZKDw+BOUOniLuEiQ/wHhVM0mYqHI7x
+9C1PSmznojpyV2AC/ZQShGBuRBpJbtEB4Jh3HbdDk+KTT7Ev9wakXjYn5cF4Bi2
kxYFdli3SRV/Fz9jzmJDJXmHz/obolVMSODGHeDDL61Vn50F91PE4Yb4cC/u0tm7
ZRqzU3jAJIYLwLimY+FLC8FWXPXlYb43Mdc+odeUwpgWrXn/DYqFcxJtUKwWI93n
VSlF+YcLSIXLFDUVAOh+l18CqOsL+rHYbrJQFqAsbhAXQtiHcpKXakkrw1AGHypB
6gxQVWT2qGqnynKFCBxOnu/NpYZ6RMjHBOI3OwkrfyvF5qhncJQUkyrgCQl0v+HS
XzIQuz9N1oX9FyY26eJzpyqoqAvocc8PU3UImKPXtcDObMpzlm3AR/sFTQB6eJ6i
l/wRw/A/agdg0XD9S6rdKjlp3imRQlw7nQ6UDMpsCnmsguxpKfJMBjDv4kJAdv0I
xAbEsPw0g9agpbGqrVfQBdjYp70UcyG2L0nKS/Far53Vcg4Fg9NNW5FXuoCFZAy8
0OicfX6iLsb04EMM6D8J4RWHAh9peN0rgQwR8O1KWiOSwgW6ZjWhNn8b2ncuJ7/C
lG71I/w1N7cvahuti09OE1+XJT3cU0tb+dchucZWkfkQG2ibipbLuYml78bXR1yg
qPb8vnz5NGucp0ekSTqVTLG3iZkvdj2NZP6mr7GUsaSqumMwtIwYQSDC9uZfXSyl
rhCwOm+Hv6OfiR4TJHpoinYhIw3LYHWGqi9gFKOlYOlzBCsAOHu//gHDKsLxZHJr
Fzf63QS+Gz+PrekvCfNz36WwaO1DCgxIjPazkHE+ARebj/N1nS389gfWWDUZa6iU
X2OuqvedHwjDSwiAQCy3n+3dYl43FPFEpgS5+o0w2X/Bbe23L6cxtMmP1RzFXA9z
faByZ/dPkuUtv2L6vujP0I9brXhaFtJQ+vmEjDWSiyyzI4N2OBNJ1fZfzaVA86ia
0YZcIYhaF9LA3M/jo5A61qE5f+yRZTGLLSnUsUH0tikJia3/XFoi/7HzWlymD6AU
imDPpEZi8s3BTl+zebsNzEyY7+aEeRHpvhzIaHROX3kJYzW47R6ZP7SYMze9i1kH
5qFu9RBsOu3vp/BsW1oTLsN/y5xlETUcUA0IfAP5H0Ukl3Zqu57EtpGe4bofGnRq
WBqYR74KHvrww9aRL2pY+KQIW1vFaWbZtvacljHREqX3R7+njiKdPdyDhZ2COCkr
udw0BW+utrSQIcDA3qCCk8ShaU8iqjfyAYziWMCsIUIpY/BSW9h0+uMr3uBMPavC
Ib1Ghtmj2yp8BB9plKX0+xflIBzqwTM1exZ+qSaBJjnB0kz8D8UzFMz1PaYJq+ov
utjIDPvsIlQr/ioFvGmBaiWK2pfWFb3oX9HnqYCPYvNJJnulcIDkbsVp5ZarPduX
RIWH2EHoNmbWZ1z7VdxzZFeH81YN/i6FGV+I6W6l4p9/e2UsY3FmEKwXFKvTuIxM
qGHit00zXJ5+tMIttYfEi6mEpUcgaTSTh/YTq6skoOTwn+eHkcPIZltpVbCoQ18q
iXxrU+mCynOj72SMevMKB1+2xCPTfh2atHJlctzBfRVm3dAPiAdFURdenDkxC6Gb
YDBT/9xZHtfXvyr3cVQQKBdMUYrCRH2vrN7FarquTdKWprg3g9jGTtRfcNnsxBtI
bMOBmTutUX5Hu+SYK5KGu+a1uigAxSxwRv/mRqQbukEM72VTrg8kzJf3hazxgVPM
BaaIs3GDMJNmSMjUrN2cS8JqdLgBS6EYOttE8LuivRCbcKEMGNsE/JdMHQ/Ur3++
Z+2s/3FEDbky20OjedaWsanEfSEXRClED+xfpXEZcFxFPhi7gkgEnu2dxjs4SkS8
yXqwjE4N1BHGnT+QbUgS+Xmf7Y9am9xPJX2UaULwkBQUhQXZdU+ie5p00/9a1jVC
PhPTrFrnZYpq6KJOQ8quMBtQ1XM25SGseV+wBdsemTqmJBlzftGVnd4SEQOW1uLF
+1cIHyFmy6kPVrOM92iUIdTIiX4HdR++FhDyxUsIg1jWP4oHh+C7kDeTh8U8+S7Q
KhRKqZUnZ7v1IVLDDWoJWVVyIHq0aKE0ZYu7QlD6PjBNlwzk5tsMXF72zeYBBRjn
m+9mOb831Shwnq4ZCZOQ0pW9plqxBGhoqxgdMkW7gpH6KhbPPCTczsZYyxgXLLrI
lhvvJtVLy2bHZGpUr753ThPOpZUEisHJfGxixBxcGanbNjJm+YFVc5nvmIruIrTD
0D6ULVvr4n4D4mB4oFfGdNroo8yzGj5aPrnyEUCHb140EKNupNivzadanbaGltwO
SvkuwyDMztxCSGRSq9/xJTaGPNOP0n9Ce/bo9Q3Ywg1oGRhi8hBff/kw5cAkfzhP
2+FwRb0SdRl6lbc2j/3CmLqcDO20TX9WCo/Y11B+pD8jeDGlL1pUwexlT9MPuk99
butpfUbIJUelsxCZeBTHZt9ydEnao0ANSAl7dYJC7ve5CniqMC++7Wb70jxPvDKT
nDL9mE3Yqdx/M1Q9VKCtp2yWEkd/HsbGVIfY2LR/rFvqFxfBEE/U5zQaWQY/gG73
eUG3mAyxIUDhaLbNpsv13GHbHXQSzRjuqINuZcKr6oE3Uk0Eub3ToNe6p1ifiG4C
5gIyL9SHzBr0ilXHXOU5qnFe4uTxWlAZL8wQQsSsvfUbe90F8K9Ad0VDUxYIpYFC
UYtEMgZnmM3M5fmzMYFYQu9/7vyi9d2zGFzrdyV2ErTqHZ+m+Rw9bqUFZoea15hn
aj40NfEKjyOtc7Ph0qQhczTq3GCKB3Q+dByMT7Hyl0C34UCJrtwkO/+fhchaq343
nc5u+17MncaqiV6Tb6Ozs1H1CTklYEAeOLfrDxHNLHfrizQ/E2OuzmpqbmsE3CCU
RYnkhFZl5NJM2hS6X4a8p6uoloI6mqzO1SScuQsnNyuyCuHEPJSBOyURDefIL0Vd
GCaCpPPFp0u3O1PwA7ebw8swhY1i25WxinKJfI4PlJrWtDCBoWtOa2R6X9ka5ZB2
O9u/YrHMIEt6t49xiL9age55Q5FTX6G8t/4ke4athIxyxtfdG4/0fIaYPO22fyYy
8PCiK/B/EsIKwZlmbBKKYHUc7Cd1GUF7125SLNdT5pZI0G3AaukqMpDAN7I7HksE
Ypy2ZXGq4u1PPPFg7jyz2b3ArbxsSJkLFm+lqBPKiOuHdvZ8jYCoeDeoS15rH8wU
PNREEkJ8gjF8tUdemWIeDC2+PAHn64MwFVb7vbK8xuR2xsI/pgV/TjRpa48Lzuv0
rMaB4CaF4BBe8WLA9Y2Qfy1BzBVTeDlFVFVZsKffuKKgpwKw29eCPN03z8b7rFty
tiDd7L+DiUKQ4SgLlLSjdfyTyoKzfitM/cDJoCXgPgCzSCAPIsmRFe9Kwp18fj0k
I7qivpOsMdRqRQYimU+46DyaMuasDT+ghsJZHOJwhEyMEc6sEt+pP0dIrT87Ggx2
vizQvET/jBnwiCJpczaQUOGhrkYem4cW3zA9PRR/GaEd80xftslp7KXXeq8HavEa
N1H8BCY+22TVJUSlQdKi+po6wiz5z7v+cy0Cqg7A+dTWosacvGLYaqXrf9Zv2A4a
3Ymjcotqctu3L5SJuy4KmlZQ0H7iOP6AMCVzlo8pQ1HD01s2wqtqmS41J6JFGy3s
NCqyuc5TBDF0DfriSbsxBhA9WrV9Fsc6JYjMBHEYUsmU0WvC7c0DrS7xPTjXOxoo
g9QCnOhRyCLu8fyJ20aJ917aEQR079Ddd9IOXjrRvqq6gOXkbns9k9+Z0ObaTTDz
yqE0IS15webwvqh4z8SDqqApVdOuxP3mmygye3HREg7o7x9yc4IV7aka65owLIwy
OAfOxBApXVhFZp0UM5ncGLKODT7Lfd8L2pzXcBdsFLZ7DAJ+fb7fxr4J4pkOkJx6
m5uB+jGqQZCUMzOa7L2unHQ54RQlBh6tq4uJVMEybhVd784UNg8AcU8ThqD2jaT8
PCUUGagU3GP1fJo0Fac6fMCQuUKZih0ZLuGa12JOR5nFr+EIE8HayZm9gJGTf0CS
wTyfOvoDAtvJbmaVHbqfYKGVEYNUCSMXroj+uSvm5o8OcAfpj2LzU6NpEYO1KvWM
nvjyASRIu0GMabSkO8/UpeHIyu1QNat9nExjjJzbU2TfjZFNjj16n1pA/51FxDDd
QxH55OkxIYXw5VrpWoKAwZYS8iQar6IpEmvvBXNWouq8+Huur+2n5hHlAZTV/qaT
h6IrexThxSbgXHPsZ05taTk1E7Cx+xfcC+neCxXCfsZ3gCnFPHzIjMjyMVyYOeED
XLtewiZFjIuNmtBlLbkdvmYzBKfpGhDBj5EvgNIRfYI4eFK9ZcgcgwgmxmS5rW8D
xXDHK7iM3sc6x50rdg9QE5Fnyda7PkyxfPpDavHbL+gA0cyDsGF8Hduyt+jzVnwr
ZwaL3Bryhs4Po8uRUHN4APrR6V1BrLmwmN1k56oys7L+N0ogzD56pPeBFtlcC/eH
AaiTBY1L/iCpGe7/GjhCynzpWlPQzZURWyLJO9Cf8fU2X51pDELEMb0IyZ3yaYzA
38iuQfV2fW76etwJqEAWJlshMNj3AAPej2VkEOwxBpvNTXlSRr5FnZGpbXS2frFj
CGgTJLYDqUMWAaBPoc/dGTnjeLgwDo2Gk/MhLbkVMN45SnC8wiSkmOqkfp9PYlVA
Z8FAtR5sOwDWG7GtcbLc1JNb+R1WJWs/1rxCWvbhWu//vMhmYUpOKNwCZzP2R5jd
EAsJBwpthIkelJY9015LgeJlRbhHlNuMgYpaSstCBaSo+SPTsaoB32FfjHnJ0vOO
ghA9MPjpZVfAYnz2IzBDHrkjZHcEZufiwXhpw2oH9jQi9B98wjotHbj/j8VH/PqG
WyEXjbjuui58Y4faUYWTa45m6L0zdYnpM6IxjzVfdaDkoTaLYG7MLkXQrLNNUdJB
+B0CmoAeVdQJ3I4bdYhFM3BOKnBBArPt4ZH8OEOAwqpzxvw6IOT1XRb/CaFd1Egt
T2ozr1YzI0tC8aXMEAN+9UrBZ1ZQv9rIfkgY3f8uQqcAIPy4Hbg9vAkHC+FPo2NM
jmSjToAwMZPrXkoNdUxQ3M+pJWcJzhT11pDMo2V6WlyAi2lf3l604t9aUsMCwubg
5rIrd3xfyytMwSPDuTBSn59n0f61o7Cm8/mvYrhOvFhVjclsZE4i4SHcZPLujtJn
yKq7KDBl9lSfj+VsG8a4Nnles7dBfbwHVn6TeI3zBQDAO3tJSBoFfdL25Xs1FtaF
g+Ap2LwU3JhM7M3md0pPxQJL/fzGyewooVjSmsDu8h3+nzg3eZIqtx5+Ztfn4pid
CBxxVHe/NjAITvGX90MZDI7wYuutpwfUdrbONYylosVwqCkZ+E2xzKpqspzQm0Nz
KE/Aj4jLsIT4cO6uglGuGHzheaiALoLpL/76az87AYijhIbXYH/brduPWBUfmf1T
5hhprnMLvfCM9sgxyiiefcrtSbQpVIka5Rl3dLUrteb4W8bvLCZe8TJlmKYodvDZ
owbbOo5MiFOgQRsluz9cpQiyy8sKe/XpQHcqW1q5Sn706pyXD+5IChVxIVqaliJG
CizGlnJ23fIP0d7iDTB0TRL3s35jDTO2VS8CLYBMEiCmKqoC1fVKeZP7d+HWyw/J
QKGqmM6eSeFTk9YLbiuUBn6buWJr1JlBsJiWw42aX9OtBhtLbjxsRU799grbVpzu
f0b5GLgXd/nad0XaFOj2w2e7eEYgy5aRkNMW4m1qno7cFZTphHd6gCaipWpvTBr3
mAA26kxkAmXi7+LfmP+IvMOkSy3MYgko0m2tZcSVaYkoON5DCKzobKTmCKqH08Vc
zS6pmrHDAVg//VRB7JJTxTjsxjtYjfTkLfFvamzI2wTFcvJPtZrKkEw/5RJuNTl5
bRNfA+CDC1ZcWPBdpO19/KRmRidph8+PIrJbl/B9GV2ppa2UxeS3TtiGkbrWTMl1
PdkOLnGTVzghAuY5rPkr5I6zb4LXzy4tCQM9zYYUJsDXWsYTtrAWvpglNF+fxi7M
//pragma protect end_data_block
//pragma protect digest_block
08V9WyL81tDBj1N5uIS8Zd5dmgE=
//pragma protect end_digest_block
//pragma protect end_protected
