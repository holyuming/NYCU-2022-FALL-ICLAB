//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
j2dfyE6T1G7i0MV2HoFb717BmtbytrbPruSVEG2N6MIUUc1JDXJhaSG6NAp+RkR7
Q5gt+ZWINq0jsZ70Sbbq6Caro8zs/YX/U3yGoSBQcT0ijI7Awpx4O98dokuAZJ8E
IRynnNPP1t2WHKclCzD7ZmYHUnMmcYPO+u2IkrQUp7GFpAuBgrOk6Mm7pFRHiHAK
uO/uaCoolRBehkMqR1fdn3LAO6EA8jv6viHcU/nBQZTxdH+NImv+SsSa/169Gpuc
yydzOugKUjN+Lqu/ce8vPV4yI9B32xB9k9bCYg89H+jSChIqDa1Sa7EeZwLZqNKh
dW5jEdqf0EQW6djr0GcL2g==
//pragma protect end_key_block
//pragma protect digest_block
HfSOmCT6lBlOWKNqhyZDD6Jpv4M=
//pragma protect end_digest_block
//pragma protect data_block
c5GkOu41Z18pev47F8c0aP8O5mq6nV72aVucN/sqmBp6+P+gnYijkOXrqonpDZUb
kV+//ahTjApFAhbNTjcZw/uNYgGWjb42tCGWfPJ3hk2NwT5XZeC/w/XP2vj1EMNa
IdJZTS7X62JuHvpcfTXTd6ZzYTXNJwjlTGXxP5bhaLTiDz8sgocPPgwkSJmIr8LM
zbFWYI1GNFiVt7B+JINX9xPaExLQGICLDzLehzN78S+t0tNwx9vJiHUkQLQLLNO6
9LJpLe9LUb9gywwmgjrMN+95YbsI/uX20Q975IHpQ9JcIZVwO1L5VCHhZOFvkC7L
Fif19Vu3b+Xx3FVKQdriiiZ2C/A7lhgs12+lB6+oTZqlZKkMqAgDIa+dMFL80ArM
6f6IJ7+/fl+Jx+y6n3RCmmY7G/mS8Rpk8OqMY8AWSmDl2wJmYVg6iNa+3TbTSLT/
m6GTXuUyVJJJ7omn4MZAAfApNQCE41v+ZO1JEGuABzJ6Xsero2kSbtiO3zQV+nWq
s5bs0b3/03G8db/9pTjaw39MTkB93tNxldQYRBd5XgA/bvHHkP7AocIMtl6CrENU
6YQVxhU5BqYEh2StNhgFnjsB88QIHxjJ60kD2fcc7pgIhbk6Gd5ntiPb4W9wk2CO
BVSCiLw13OvyDLqUQqXxeTLB5oxjLKKb1VUjODk2Rx8EX+wVH9F5rbGOwVJmpN3J
l7J36iWK/jAuoUkuK9a/TxwMdj7WgDqf8tK3BVX/zlvBfoKikKRlYGRxFxfajn+K
OteLMOkuppVbgSxJGxS9NAcSv6VV9Kembjit3Ff3A/x+c/c86Mej2jg+AI9Pbrfd
6SfyITdCrShI2HgaDknYZ3n413wrcklOgiRH9Qqzl6WvKIocaOuDVsrbMtuqjZY+
n2kV8ad6hOOTG+KnmHZ5TuEydkpcC88uDOGInSivxbrdiXIaXS8sBGYYrawt4o2H
7a6LVxcaje97R7ceJe+4Gfw5FZlLNGnv5MZ3R1jhDzAEjryJj4XqZFRYSeZ2D5AN
yadkExQGwZ0frcxtUYMKEb7JpUTE12hckv5kDK08B0tz20AXs61oCBRsmcXfh3iy
AnnzaYIEmhJYFWIUjk+mhOGZwnHCrf3XK0bR3mDU+n+zx7oUzwMz1kOc1qe5oV9D
AzeK5/3gFMIpfYT7bdtwYlebbNes1rtMbUj+4Z+fD9HacLERW/oHt5xir92a5fKb
82b/uAyGQkrEhqM/QnAS4ipISHep9NULMimdMX8MvIA8aIgxwi5CE2gF6yG1Pdki
2s4ZQWMMu06UvkJXpyst6j7wIg+XolZriSrtqGdIJN8cdjRIR4us5iaRhyr0pAOD
H5Sul/+VzhEP3tDl7r2FILEfyFLbvQjhywaNg8+uRLdQK0piETOhWA8TX7ldu2tY
AZYf4jbW7fTfik6x3fwIWh2VO+LiqWeSD62s1YdvZrHBJomE2Gzqz8+jjIqSniDS
Ms68r4xZEdXXTW6vrF8y9F1S1gcRJfEqLY8wTJIYj9HB14JeEfCnxuwbr+KSwlq5
bE2xqEGq0SNzcuhgZbC1RAOj3KWOWz0QepOEXnT4B2sbOuDYp4ZZQuBbeOMizA+v
1T4Nd+ykynLAq8HReSVM7l6lyXA8J5Lz2kYf02KpyLXcpiqkSCQk8IbtWwcVA7gc
ceasi8heD2pIEe0IJYon4jPzvipn0/zw4Zl2S/iDQmf8vVKGOgHPq3ec98GkbOZd
70jAkDX8KKvblKyIDb/QVm+dVrFa+IFrjLQPEmmHPY/J1XMtvDN3C9+M/2jg9sDx
xNRH0oaBStUw7wLcIIcdHH2HAQd2H7maGGlt1afUiMe+LNjk2lIttmQJvD4xGKZv
ifjPXDK+pzemJuPUzvOOxS21tDk18n3UHhKdAICQQzaXKYX/GHSmnaUxpKHVm8aG
G1zYpgWHW2nxY4QFBuW5DehM8k/Dv61qLMVPmvhpGHoOyFKBOCxiiQpI67cD1h8A
kt8IJCOVXP93m4Y21zZjTv5bMatHiwhsX8rq9kXr1uAAxgf3nuDMmWJXjkJzkJ1G
vZFMOuKxX797lCZPSpjzKzbrhsQo4AcswfznzcMWiPPeXS/AM7l2NNUtXSlU5Bpc
GeqLraxY6/0sde1xH2myDii4Ros13Y7VmJ40GAElndMpBhyRRquIIy48QK2gle9d
qWjXVRjkvJKdhFlMzdW/O16mvXSQRP056NfggN8+FlTvqvCoB2G5SPEk1TM5Z0hD
DUrXd3Qngt2IjQxoXK/TOTB8CBT3ugi+BWDPSSdEG6Hs7GAC5eL3HN5BvA0eHoJ9
alZCW/g/p/VrXjv9kxbMwYI4hxE2k2xzEtJiIUpmbJFFAUYQ9HSmActLJqSxyyZ6
mWWTq2UCUg7sogIMIDgAb/wKqPzIm5CWEtlcuGb8Gq2yuuc/ESZetYayzye6gRUz
Mnp+QEkzI4M6XWRCc1KBNEfttwvBxYV1Q1wEI/IbM8XX4oxbts+xgGaxx6rLefKV
g9j/MSCIWkoTsz37BMdyvk4C/8FS2y2/dA18twGwbATBOdTHi+r8otc7RZ7epF9W
EtBCTccU0Tb/ezMQSj8cy+LcJbSLxjqE7OGH0tNDzWcABKFS1WPC+QMOMvsd0Ca9
yYBl2xA6f+TBALSRSFWo7rJW0teVIf06psbVuC+vn3q1hvdmilceBjbgyU+MMWkQ
bUpKUOE3gbFKSHHwCWojqyXHilW2T7uGzqX2RJzCn7Pe2VhXWAjUgF714/m2td9f
wSQiryAieIbgbLFHvs84GIFWr7sJdUvVoht5xFfkq+8B+LG9PlopmXAbQ01VlJHu
JAV7h87DDIAKVsrRX6sIKivdV4RJGn/K4L/flXmQ+jVXvPzRP11/lVMITn0FyewS
fhuMsIgFMlq8CXsfmhJUy/PRN0ox+0yEdspRV3dG0HG67Kf7Mu3PgnizUwKJTDOp
tZOT+2NByxIOYlBHigxjofu1MIkv2/fTvrzGqO9h77IpVrpZNnsgDJWvINlpMttO
l6uC1QM0jLHZFaEThC+IG8lspeZuzVPsl3QcxWt1ReUqzX2j8VrM7pLDnch84H6m
j9wn/cJbs+T7GGzXC9oKNxPlXTaMz+VAitrN+z0/zoJk6nwQ75Onweov7g5cZZ/t
Judfdy87Ab8NRbrzjxybpFQJy3mqxx5qnNFeoswJj3TXAhMIgL1jNEKdNc9qwaOI
6yICW3D0wywUyvARO39zUng1zdK7SxB+q64OLc/x/xmUOOR+cvjwCrLT4oebaBBF
VTu9RGlS31yk83RfVNlG3gODNzxfAUr3TbqGTgasZRZ9YZrV3FAscjE8oj8CuM10
4UtniatroG1IXnyNt+xHh4Ge3Ta6qyN9zDP5HLbplz3OZAK2ENyrHtia3Qx1mws9
VbgMB13HSkMU/Y+n7Vnwv6e6jkM20XTPmi+Ery/mbECnl668lgebIWCDHXFqzn6I
BoAAxOb8gXRrfoU2zGSkfjWxRBq+VHoJXHQ/3V2x9/OpMAOzpgbPAwR+PADuuxoY
5QBQTa+8tRmnNJ6ryxAXaMv/wCHRt+9Eg9MSChNzDKEI0X3lwA2KAW+JsMfUiqoY
37/4j9jjnNyGgrdiWQh5FPZEF2BaxP6sszhVGnPoJVDN6y0iVSl3GCC3/89eSpxv
kgv0A1IRH9gW6XOeU6YPViXDTvkw6r4e1yhqQzOF4GErt6s9enV1tiGuq6lAMTo2
QDD5IpAlgTkHJhkebbuTFHnRBAE9n93se+LIIZlIGJh77PNp/85OkCJs/ZQIeWP5
hJbgUp/QyTCvgRa20GlBLCsMOn/KZaTMuyvESczz7u1vhnSJHfTxdpb3eaM7vhN5
o5bcP/zBZZdQU1vy90Ll8N0MxNzxxobhqKpX8+lFT1d9arFUw3Ye/zGmb19BknUB
bNICDCYtA/T2mzp671+W7MPsiaG2HbPXo2x/2prvHHwSQ6BQhbLfOm8q9D31U5fI
bWQzsI+pJyZvHEq/tAet6mj+PbLxKlzbqP0vndDUgx3getWTHqKLzZCzG7bk12Fq
kCs3/h9QNPb0VIdTqdeoF5J7JhoMyBO7WKyD5RrsY7Z2cd4EjAOqty3MlY0YGAI3
w5xZ962gG1CDoF+DrNtgCwGYnS705ax4plg3h2Y6n9kLM7usje0kEtqqibA1E3sS
Fx23gJmrk/aG7VwC5xrsZhA0rRDDjRPgCJ6JQ9JtU9yOFJ8Ni5YRu44bM/gZ6fBM
QqwvT3q7XzH4deh7LocL0FmMPZstTHaAQljqFQ2yFPLtbaP8DxpUbrF6JjGTjQyp
YGpW68Yq3BCEh+nIZj5Nk2tbyUrNGkAGH51qP9LnY0MKyqH2jP/OkBTwon+vWhuk
O3WlKmBH/At0aU+gAVeyPtRe8xyC16mvX4iS+OZkZe9MrfHpO7gl4wxO+l0zwP4x
2zs/dsYu6va4tAI4OkR82kGCPNf2th8zlmrdJsn4Q2tLve8SAs+Evm7pLal9f+Qw
pToqCJJkoa02s8wG8tOH0dD4oJlDEAVvFD30Iluq2aUTej5TgPPKdeNwQkKswaBO
zI51HBQCxHb5f0g6pbVoLkXo/N1ae4/M1SplQFGGfuYNEBAZn4XXopTQ2+yREO/K
1brfF2PSxf84hBDUa9XcknTHstbN0mxtm6cqoCdyL3E6NqLZU2ck7+jmyGeZFfw5
4KtoSnzR1sGG5wi8d8q6T7zH9UpDqBc03MhdzUYiT9WQJhX9CDuWilEdw0tZMjE6
9LGBtH51ELWc81o9O1x61MMn0donerQssCKMxUZWXIuwYy8XUm7eXfnVVKi9xDNy
234+MzMPHr3C3MGYdy9bFnBMX4HZmIOQ0o4PNM+pBhQ1DBaPygGTlZW//P+ZVBDV
SSq2ccrEZEzUM4F+adykNJkNczgzO+KRCo28AXdRTEidbGfQPMehPgyFp+c7bgTU
JA+NlVTXs5kdhEdvvp4kXDwetbwGxXPiVddUG4OjEr1CrzcgFuSInujnnw3MIMzF
T09v/8CoJ+GnUzilScvThsmukK3LmWPaJ0yLzItx7jE85HsgN8624Hj0ZUL9UwRk
8J7fgB0D99fOcVFzfiqkf1KNJteaaao5/8k7VrXi5EopaIVUQO2hA9eg0clFeWqB
buVKrbwHPFbPGJoOMmBeO8mFE9gftKJ9qPvuAXexYN/xMD1P25kLZmDvVrhPr5UO
NVyAzPUbfCPJMu/e/oX8QspqEYz+Y0tQwES335bfD0NWLoD581r+xilBhYTVKXPW
zRb1aNTiK3Bflz9zYloQoG5TBmPebPt3Q/8SPRy9E6xiLl6bYQpqpa4J7ldWc2Tu
78p+FC9Uq6n1eiBBYfQ5viuYf3oVQa0zPRXHsjwWZZPhGxR07F9qMFxmBp9E3lni
xWXVHnuGVjbQBfozINPrX88gKOM8+mUmH36oaXfF801e0pyynSMum3Kmd9cVctt7
15z/zMJDoEFrlULU1/E2aVM73nL2xKo4VgebODPEsaD0FMLLI1X+bOu1u2RfvOoe
T6mYJubFDS2rA7l9+hIj6pBWirPq8zT8EUopLVvD4qpqlJ0BhPuW0m44aZDdHVME
RnrTELz640ivgKSUa7+lCkArltC6eaEBTCoMDoDdtOORIhtmJJGGAK+QPrfiVrpd
ikUGa4YFBjh33TWy5A8Y+pclnqEOYENujucOsE/W4yYju0uTDGGHES+0VD037RUV
jv8QYEcIyXvKfVR88nXoCIvXXZXn91uk8wDqGf507rCHzSksdz3meayQkmh7dOXq
2AMVRwlg1mC/Rtq5ubEkauallSoxsz4F/8GC6rSeoxKpS/kj4odaKWxHh31h5kS3
rLDHGN3yRCRqX9FYUXEX7VTGwOpudiq57l5ONfzJeGVavLXIywBkqGfj/YL987BB
99QiRwNEJNcuUzl4+Tf27ebJyaZYiMxrs3H1xRK6wHs773Wfv58j+znF/mzhXPw8
SuFzvNqVJtDQOzNDLBCLMdu/kirGD1J5pYAxV5wTggyPeJDuOUZkY82omDwCNfAd
G39DCV8YIO+qdykChyb69MEupcT8/K+BfIqbJS/XNXXNRsZ8IRtRxl9rrjgcMj1+
dBoiz1k8Vuyhpfkm2yuZVMNVXYyiA9WoD5610GyvBaY0o6MNl6aP0vSyxPJjrqOD
t/vBTq5HZ7RCNH977zMcHcNwFy01YhS0bJf/KTuW0dOp/Kdd1R1V9g62bfBj+jvI
Z9LHzVCZbuBpJT3OycvLt0IMPE45KO3FMv/xLPIlEWbutb474DvYaGZD4PcG64UU
aDPyHrxlYo4fxWuNmMGJmOa8Sw7HM/Iv1oRfncB9FKOVMcT6zAVV3Ukbh+tZOv6M
3EEyDM9Ar08QA6p+QsxOKTK7u9XwX/GPdwdO7AK1a64MM6D4r37FW99DOlvsEqLc
k7WbGkyBt0Puwk6iTNSYE0EzZeqdPJwRZUYeTbQfAqOzy8wpIOaL/a2PyRxvuOhG
jS2U55rU/qtwZhRQ8jOMeZKXjjIcvX5bDQ8TZXYhzcOBQ0sluzpphhUjwW1PCAPQ
D1Mfy5S80L06Pgiq8RVE4LHv1GJZdUiOnzoKEN8PyS12HrrHJiPI9qvPL130jQCO
PKbuiOE4o7Ph06kI0D0KUBnbi33g8hnW6l9YpJxQBokLoDmomzvJDFhRie/rOK/w
nBMcwJCYLg6tE32Is7BKBCX283Vr6yisd5XZWZ7NSavu0z8nX3M1HvjAnA/nKJFL
oYcOoQoKJKP/5YEqq4pv7QYWR61lq/WT97H22FKsbWjdGqSQDA252affiN1p9T/0
k+1y0NWvHiWt441NkDnPWcRxYABAKndsVU6OItYmdAmQyxCtYvF3gbngs5vk/GDL
p6LkB687tqQeE/0D9ciUm9LrokBD3cs1PnWKGdm+zWxEzwfp/zLd7onNeVo4OMnC
T4h9fSnHsYW3csmtBY9jLxyLpFExG6xc7meKvUMoBh3reren+icTv6fMKQ8SGMcI
vXBT8G6D3FoXTW0ZAr8BbbVCIgZyqRcq6xyojPeV0smw5Sr55V+clSX+REsM/dsp
Q4qRy6P1dqI2fvtoVXueF9cQdaqr46x4/ORBs37vR6P7nXuyFMheRqOhE0HcjWsF
vKRcsl8g8uljVfpNKMHQcy9xmIXEziHfLTnzNFj2R2awo36LT484j8qWh8MOLRqf
pD8rQLsxrDIAucuxQ2z/eGSmjl84irxLxCmSd4Xv4BIqwAVJ1nEZX7SJNJ8VIDBn
imefqaHo5qPyepDhiM1/lAG9janiQKqsg8FtN3IlUi9SztWNN20c7hPxOY1ryqqs
LbheWGmiWSTQPlu/XupsqCi6VSoBE5jgzaBHk+h9Yd+wt+y2Y446Gokes8hkUgGl
ymLTxNm1Cl8wfklf3EpT8h1D4GLAfzXCnB1G5vc+lcenwxQ0YkdJ2dtNEHx9oaHd
3KLgAoGU2NyHTs6Cw6j1f9vcbh5dduCgQN+aJ7Mt5lLXI6oIxubcAicpihnHNKX3
Ens6yuycEBdPuq4JjZvvnchn3QcSkM8+vcTS0DKHvvbk2g42m54HA2E/CXs3b9O3
t2VFHhf4Nq43b/3HZcGA5ekGU8C9JmTv3ufzD6olroxp3FpMxwOK5hDJ5h2YTiJY
aqTp/Ed10UoCMIOX17+U56Y/5hG34sGm/lGQ4Usw7hbz+hMcYQsxy67IIXKNnffC
omOBD7UXtPGqoFn0CNQbio0PV5E2VxQzS4yr13ffLB66JY2qEBfFfFveUZdUGJ+G
/sVfh8Zz48rVAXfRECpa1dSyANgjDzNSg48NQ6xUZeRXiFhW4KUS6EtNT35Ph6Ww
zz+ht7D8zh1xedsscQlysQ2Uo2oV9Hs7IQLzL1rmHGMDEvARVLzsdac38oVMS9Kk
44XiSa5bGRH/5XjBogGdm4OQ/6y24O/90EvTYbaWzU4P5638AHXl18k1ekkkGFE2
wB9AAIuPLdh9k+ajYbm80nl/czUBmPwt+/7BOS/cNsoElgIIi70Y/xrnDR7Sc4au
nZNpL5znSPNVJ6LEH1cmDbKWz8gucW0DwIvb6QVo9kF/iEDCxTGUJ9aSg9d0d1A0
LfcQj5793rDYOhK8zZQOTkGz5c2mAL+B5XKX+j2K1Crt2agCQhqx38g3dPyJrrse
YWR1prf+I7LxPAaBiCy/8g3TBY98uU/Qc12xUHtLsEk0rggYJBuDADZefGvOI/CE
L4tb6XFM2NJrBiG9Qtt5rartNo1NsArK8lIC+vVmEwM7zIT2u2+/J52iqb0oQg2M
Fe71W527G5C2G9zYVkwLKg0VTub/yL4TNeEHoBS4bPW2JVS9UHPPs1gMkU0vpGWb
NaDlsOTT391LtIoTgzRA9ei8TAE4qnmM7dTlqrgn51atxD0FCsQHEInPoIl5I89/
CXcxmmyZT39nEDR/Ib6IE6UziyhAnNaTyZiwqH3xwQqSHUpyzwabz9T9AobT1Abb
E1A3wSHgeYdNTar0Uz3LTyPqB5GHo8lG9nOZpvi/3cAWveRaIYeHmMFBdUqGi7se
/gHx8fPPbxLLkbBeAVTnROuZS/nfWt8RX2r39xeiMZIGGjh7aWYjr4MDX6YftjZ5
tWXwYCa24vJTZPE4qRDxGvi2cTYsAxldYctsQWUkdpZiCbe2yJ419snb09sGoWSx
8Rg9u75RrUo0hkkPPVjhEC56fMhdCudS2w6Y6d8nY8SqZFcCmD984rBW5KRwAmPi
hW2AbSM7ijpwZW5tKMuTFRDVMgnzcggk+VGen1tzxDqOWPa4waTqyiJwW+6grnhA
028wDajN+4wLxlQXEcY5qg9k41HPPvx+BEh7CBLByY130mJ2EVHR7nscpOpDo5Ud
Byn20Pe/zKQQ8+Gh5LdDko+bH13GE2nvlSzocW94W6c7NdsAq0rYD6ea/+JA75GL
1vPd2fECDAcwhOYr4oZ4sxLCHL7G20reSiFyluyUHb3YjOnkmBHyTNwHA2R4M5Vc
Kr3shJqf3r0Ffz1lPt29RMKZTlUr0XxGcGBCPHdTQkIng2VJzgbNRn9+GTNW605i
cNGaLKgVnaa/GZoOnHavjqdZs/4C+CLeG43Ar5FiFPfOhg1d64zbm87Ycffqzc2p
RBi1jTyjJ+1ceeMqyPPUao+lDiJVk8eEcHIR0BlvOzb7Q1Xw1geniQyCWO2pia/4
zcCdwRNMg+MLwFSpObh4zaZ+T/3yYPCww2vexOBPa3ShFV58mHgFD1NLz/7N+AzO
n7NB4BjHZYFWteoj8JPo0Mij/puH2Vg5lA2Io20uSNj0WlYMTZxB13t0aC3g/FHm
KOzKjmennYPX0GPzeSHjDc14rwv4opkPYzWCKKAAaLBtKRL8CqDevYPRsH7WuFYE
hvkr42TEhpUc3CR9BcyvrHeM1FeNYDv7oExaEFtaxDPtQwOexBA7PjY5/NkcdSV+
luWNM6FBmAyMcn7tW17hEbmlTDVPNae4YTiJmBqGtVW5nslUqo+XCYtVpmPZVzgc
XmM9/AjuFh5eiftQoPiwvB87nLujsti/mHJOulBL17FqSHPRtH7YG0VHaj5x5q1N
fLHdgktlLkB+IDJeRZSmk/H/b4KtjBDf0fv69wk0CxrHveC4a9dWNuSz8i/CIkMv
icLiOIxsGAFJ0+S4ZdDs2z/MHICw7vOzCw3J26g+w1L8b5KS1nKax8raUPY3PDUW
KS63Cmp0tVwTv+kJy7bAFQK3M38UDhTiwoz6hgi5OOrXzCC5v9qAMfvemYTEfGEh
EYgM18qKoSzd5IICLhDcM1e7e4+iP301DtQi6QvUvo2e2s329rZY4tBIkqcQBR9P
KJ4POtCvb/RTikKqPY6toZw/FeTxiIkUVe76N/5VV5/0WKMP04y5I7BSzE0G8QMB
fTsHxqV9fZEOARLnhkKyE393hdu238US4hAnUfvgZs2ovm/T25dni4ll8GxXHdC9
Y+gLMVPI44j47VkNOcXK2pNDXQF9/wQejDYdi6+AZkDqS0wI0Jeps1y/VRYQvQQL
KHi0sN5i9xVTceyutZJ5Oo2TeGVVvH4pHhyrhsaE3GvWICj99nZeJW/6mSTKV5so
ayMbiDHvyS1cI4+cqkKQLsFfgah7PeToROIPXOFHLSeq7qRQ9Y3xKmOJd3Rd7Z/d
VZ8gh+L7HAB7pwTwd0ezutpIE06oSYlypoxsDQQOV2E3DCcQaCvSkSXCXF9T6f8o
Ehbe4v/Vz4ThJnBSSva+NOuHxA54SBYKwUiC2USEuXo3XJoniVgTPFpoMh7fKX2I
5+fPE+Peis+FTSIzwZDG6p+bOEe7BVVHvft7rNQj8dQ0Z7Zy5Xe2H7IHRD+ZupNU
BklAU9f/55oF63k0Fzu/6TpglRIydzCJPDFDDZU+pXgNTHIvDlrqVRBDpaELZpdF
FfyFAC9t3WV7hfvjCUNLJNVecLS4i5YjnRWn6tKtCKqg2kssEcbOiCzPCX7hqNaR
4kaBWlvLDek+i+YB5//65kRzeR0kKo6yZTHfNtqam9/0maRDldfRFxUacCx2IJrZ
wsCMXAP14JAXAnfYg5M5zkJi3ldQDQlPWjFh0re7gdcdDbapVd/p/ebq5AK/wHsT
JgMtpDpSeIcza/Yl8Ckts62e+P3HYZUFzJvHIjEVbEKndqOMkWWJs42Dn4zLBQYj
GBopxiigqaNQ6ozgiJEF+KUX2okqEHvZ22bj61ZuyEDC/Y7CPkuS5+xxuwxKX4Hm
+fg5IR+Vx1326ebZxxD3qU1b2y9fhKLLq56vPYecg4tScC2d1cZmCPuh5EQOTKAD
pqaLanAwsUAw2hO8KXBEubype16Gq0+ZnTnPuveulnecUkuNT6smuvL5kOJlV0LV
hxjw24oyf5uLLrx0qPBgdVV1UewcOSxYeQQ9KvCglNAh5S7CaMSx74/pJRDoprGC
UY0QHqJtFeNWgFcH27pdUKjNdv5lpOtkCOZIBRDegUxA5sjyumibNH3K+fIEmSJi
3bIJbz/er8s+FCcDM0NYf7BlAYNJqQdgzpoYl+a7SrGQ3r+2k/+yAU8mw7jkrTTS
sGRDsDjNQZxNDjy+KrCeB1WR5IGWa7NRQYq16cubfDR9s2+Ge0naq5TXC23ZEQJS
GONQDV7WHJ0SUMSr7Aq22+oI9O+upT0DfvaAwpMqvs98ZqBZOJ7KQfy+61DC6QtK
CL70CzHhuJwkKeXU521sllPPJyUYOaS9tfLujhJ81EjkH6qxVArgrxrFKX9i/NoS
VmC8AzDrmka3N6nBYxW15IqGI+10Ybr+lAzFvOYozgFsPM/f4E1CsFZ2RYFgOFcC
TiFT6O6mt4bOOo8ft7465OGOqsxNUAj1sF5FJ+B5yyLFDxN3dGBQCvGv5qZ/c86J
JIDgT44Z3S7QG8udMtba00Mt/q374ZHsGQnna45y5TCAHjp4wAiuA7bEEUOZeMFr
BUcJlCGeqzpbKetqyXqnbh2lrYFqz4AOoWXrAuuIuicZhd5Lu9buU0v0463EMU06
eP83ENdqJQCLYoNK/A8noeJ7HQ+k2bmdLB3Ff8pv+BPedmyzydNTARzbM+idsq7w
miITBcUNTHOZrBM7iIU0pyYXxGz9Gu4KT2JPgTbVTamQ6GKINp+2JT2eoWPb8t7Y
bBtrTgJERFiFxN5N6PTTJ5Dax0EjJB9PVMJ/FULyKRaVL1XxlE/tDvBNapINBOH2
L5cH83qukFVPMg/iivz67Ib5dqNErsuZlB4FwHvsAY+ln8uS7SoMw0zKfaqVgVsI
yRXc1Hdeq9BgTBW0RhT8WobZnVq1OqKCNpwoOK5F6/w/tW9tmcPdeGKrptFEX0vs
nRGJBiNLYJCQVSPdiGXpNS6MFRbhgFwaVHvRKvWfU5zjX1jlKNDT018ojQlEz1qB
7cAXqvMiz17GUykBzkHhdsZa7ZlIN+ggk8Ob3EL8Y4DaIxvXdVk4xZk+iLjY/oMW
lLLGrOTMLGQOJ2dHDGt53HmadDbvfXxgISZqoduPKxTmqhzAMWXYtWR3aoyW7Xky
m46ZN2KEx8YDYhZt4lcBEpZNm/hK6uPWsjiiD+96u20Z7e2FPrMzcy6/jM5uuhIx
kSuaAEyCEmlWLZOPFb3Detj4flAPkxb5IsN1GdFKBwdwUCdzGNvpHLKfuu4zxhtr
neleajvkHIUseBOd4yh8ovp9N3QO4LYmVOKSzGGMQgnWl4T/Bzth9h3G+FQ5ZvqM
8O9mxaaqr4K/l1IalhCCNZtB3yIVzMi091UsxJu1/TlQqH0qb9zWWk5aqtkB/75e
cJih4IJm8zsk93/UtAS1RntAErjBnZlWiPcb/ZwDHvXNNkJ8+r04OFe8f7YvN2iR
qNW47gEzlUIrrT6/osbfGskxZGkGA/GMN2u+MP9S7h0OyBrsv8QrNXr5LPrjzW3X
DzQFE73foHN9/J2WvGvqIABOVqYGQ8+wcx4Rm4fGR3qBTTOesGda9C57zm1FHdyO
f+8sYULYTkoQgjsE+AlTbnw6auqFSb6JYaMpY5Zk7K75G3/zOwwjNYBM39AWfdyr
Z8oacw+Jb/AInKZda0xkui8b759zAjj1liJL0xj2JBrvn+SH0vP7xSycWgl9PeN+
eKTcWPdYqRHbDUESYxCOEv0ATLliUIY+0HfzhhEE3+HkQf0+ANDPccaaCbmCcxEm
5ymlQ7pDHP5mDUgNixVuGyficTuQ0xBQ49fACGZ46Tk+p6uHpWS4U8cvVTn4jZrp
mfuA15Q7uF4su9nZ4ox9oGtmEBkaPFm9QTaYuOLIw0VkwZjBs7fX0cBaT98gINLx
Z5GAOxox2qW8k5Q3NQ6p8gHfhzGUOZKiz4Is66lz8OFlXHZ0zvOF3X7wxQeKRn6x
kkdLDmtOS/Bsy7V8vYO6ZX9iXhn0nQjj+F0IF4SGBUlLIJMUJfRe38HD4lS3qCcK
P3HgEv+y6Ay+1S1mRmbdLFaVCDEtex6ZQ3pwmCbw5zUGYFoz3+9BLuum87jamy6G
AmzWj16pBw+Pu+X7C8EK9ijTSmqIe5BP6snKW+vKw21Kb9YBr4HqbxHPzEj/Sdry
QliQ03rxdMetIy3CizLijcv5xX63FpMeYfPHvCLPcnZMQ3j51/Sk1ENv3awqUHZI
rPm80v0qxANnBcdGCcO5NUwKOtqdgoWl8YCav2iTYAm2cj67QMHfVcVKjg18Exzg
Buu+9E1FXIyEq8uioU2m72GZToF74aavc2RS51+pRf2kz6Wbdn+EsBFylxQt5MtB
y5j3EHAF+TaV4LkQ37Rl9Kzk5g7lFjhl+/qJi5kOEg1bND376l4IgCCEci75N/pp
Hvn9giqn1u39Nx6slCpTRCAeial0Js7xb0QumH5+rhcglfjuev0Cu7pUTpcBeuLX
gcYMxyZp1zFsp4LtTRThb1NENPRBH7ZEXODCdUB1viAEtmoVlSGC6L3CxxvSKbUj
KzqpdNqnr1MwhwyhDxxZfYNxJ925NXHwo7ht1sC2CTgFbOnt5kElNYw3n15vsqyn
NUDCbMkQF95d2WEi9Qi2dxY2pM0X5MEEuHpbzQcikmnt2BY0W0uFJlA59Yk8Oy/V
pbvuyItq5JPSq1OKUc2uQnJjV/mWCdiSyiV3nzJHcgTF5ZBJzxLTxqVPP2nqFBei
05lMul4OG4VYOxJjnyUQWEfQtIipOvq+l00PcKvhGIsfVJCN6AhQeU/arHcgLTjV
pGRzzKR0GBzYBhssRTlnBzEdEHKiV0AHxgnx+L8dlifYqk6LEhopDo0aEZtyiwi5
SbcF3G7YjutJtcWNuE5FRsCTdQmrWOiC+hz/4Clp5zTSnYDHNBYmtFzAAFnvN5RQ
vYBrOKYsSbPf958szQnqQNKs6+5yVRV2iw8Rfx2K3U8qR6LTMhnnDGnJqWKo2R1Q
KUZt/M+heuQDANeqJQL9ahSuUeRFki72+1/zB2IRO6NzDQ1IXXsJUFesE6CK6O85
ordVCG9D0vbUWLcY+W2ZwErb25IqHPHPvAThFu0fuA1fcqfJQ6y/0SVQndvk/z/c
rZeYtyvl/Abjb6jrWwZxNmWkjfu9vzSxZGYHutnJgtEnyDGFBcoIhLveDxkHONF7
zVHddMkm+vUN0JlcPL4iLH+R8jgvBl521cz6//+8U2UsLH1h1lsHR1gJL1Ei3OtG
iVOy0r99qBlqfb6B4anGjoBrDwvx7CC2S04RInxUD3ib3oiIE3k80qa65Da5/RP5
Pq4LxD9aBm8sA41mafC+8V0TvI9UEGU5wcWnAmgFeLRlkQ357LSdfSV641shYYYT
84Aq9ytrirAwTuXiugWiJQgiShPz2yPiPaIdVy7/+Lm8dPNhYNhE/qQdjpnv9o3F
k1QntCb6wotdZN8fLjaMIohTukDHhwDjChVlUWQAYW0IbyB6Z0+g3toqyY5clAz2
9vxCBuKB8pbULFRFHdUHkX8FRYsCyXwJ9Du7Zhf6kbK8KiBDF4UJtj+MqSurevit
FrmY6GLlhxzfro2LeUSt7R6MiBytwK6HrqS1XrKjkJI746X5HGu0lYzpih9i0ypz
eKZJ4kWwF5cj9W15pHUV8wQvQC3eqf8ROwMQGG4jJ5sCFTN1CY+kn8MIT1V3y6Js
cI4O/zwFCSP9WOgG84xhHmjYfrws3xANNpG2nkiBy6g9uby2n1a93maPcg1BE5S7
gDY3AhY29UElE9vUIBy/sVB+8EBuHNgyYnURjkpfP8TXx5qp7f1ORlul8BqCZNZ0
AByVu7KOu+Imo18NMvAzuYQ3QnF+8iMvv8dxD33M6ba57FYbT0Vrsrgayl5ppojc
Olg31NVd4ceuW6iKL19LVs7MnGlFNEN2A086+1sXatMgxnm8dt31n9FOliyQQBIS
CAVhETnx6RmdgVYdi3YNU1x2vT7xW4V7mTPznuVkc8oq3p4CUfJrNZ7epZLf9yM+
KTSs3/hfVbH/NI7VPbU28mE2kQJ7OV8ZUPL3eFlj3XefXiHdSkWr8FWSgPP+Br8a
JAA/NRhuGO3sqSrd9xubzTjv24XHTCfZLIvB9g1gnZqPzDuPk6LW5mDq5AJEVLoY
yjj9Ng0Mg75fjXYUQlprnD2S8qZK51q7nVC0LNruL1VZmHq00/y1OwavviiWhCDR
l23/f1SgpL7kRUQo2Y8Amv8cyY7Xwc7+RSnv46L+zPGf4BmC4UnqGj8JGYXevJET
4ltDJ/AoJBUBNyh0x1lbaqMJzOdoyBIgGYODEwHaea+Ll+WWjmHWynUXtgIu0jre
TwliGmvUCE+sMazhnfq/R4oE9pIvUwBuD1TjPRkYfMIQnKYdY76EM1cH6igsARqd
GvoswDaZGDlVZAAqSkDdjbey/I1w+7RpHyLC07A4fZGCRJX0SPZ8dEWQCysdIl2+
k/6rfBYooAPNq/w3h7xpNjxQFfjulgfp+PYNTu6fuwty7eMOjRFcSgcXU7IamZGy
lZVYVzXECsdJ9/ivvlWy8yClF7LsXbPi2iNJz0cCXy+hpqm/a6t76ps3lzW4B/KG
o2cCpuMCQpnQmcHeswb6P7/TV6socq3AP2eUbiXrsMHyExbWgqjMXlFDys3NmY8v
46tLOJhQZ7sh/DHf/HXWxXBY/m0P0zCT72j/DKgENmsZfy5XL7T0MkqxT3L7dWk/
Ihf6nvu4NiTXluwFUqNyqoLQNsrF9teMra3kA2dTmejfZIhpQuQePqAENnNUQSIZ
GvaNDxo8O3NCGz5DGF3VZkznQQeAXEcuAfFE1s4A4/AYSrAMgG1/UTrEIdKFNCFK
5nr/kfwTMgOFC5s8ZOPHa1fY/m6UBo6z25YSHRf6OeX5mbdy2QEcGyyeSkHdKmoT
UR6n9QePOFOjri1eNpATeI2xd3TyKqG5oxhk+7nQhZok4mImF+VEo0WgZQTiyPUN
aDHukxxcZnh9zYdHL9KIi4FV9iu+PLm/UN2hljlwaM3zuHYIdIG2JJhNukQz7OoQ
1tKuOD/X0abR2kYm3Lrlhl35Qtj3BU4SsnF+EoKGuzLJibjHtV6/hDiChEoyV0AM
6q/E46szV1US/43pZke31vvsiLTjMeNr0d+2qEDUoo3N812TAuyDGA/oZT+Lh2Zd
M5DZ/Zet4piyA3wUPNyRFkpSnwnGDVZ68vXtXR6u+BQ0a9PASF8CaAriBfkSWobt
XsGFn2QJFKsfj2wkBnlzAq5N4tx1WzGeIDuQB9DqeGzIiSCTxicyNlh6AwHVgfVz
gCHRCvhPw+2yK9Pdn0Jf1SRyEQLKMHwviyGdf6X/FBI7RG6YLTHfa4XX5iyKRTGR
G9nf71r0tKokbJjHKl+NF1sMCxXk5bEjf++b8h9xgSam2ARC/KG6zAPgVsNBCHbt
M9mRqdlbwXlBogQOKr5/8MWKiplUnDY+mO8uTbEAg4O5eqb5GqmH6X8T3QrlcVPQ
lWLAbkqTLJlS1YgZEaJWTgNpLu6kKMvmhddLXLWgJlLz3wkialUxYtuhM+T4wmKf
yFDxdAY+PostKx7qI9ciU4q6pzXdgj3vQ+KsR4qKH8sSRrNU4rhYc+UQwMYj1uNh
Dg6USzCBkcN7mD8jePLR/jOqTHr6/590gXZYisEnxPXEPGg7HNLd5rBmoa1DivXZ
s155D4FbsbdMOJ76yKHmRN0syUWKTpoV3bbqORXEMWRcxYKfJG3fAI8z+1XEUz/k
DJXalBCpX/8gj16Nr3nUV4pEbfzcb1bcADoz+iNphOm+iGLFuMUL3cVPGtUvlaP4
eGe5jUEedj2dvP0nReNgcn7U43widQx4YKPElEmq+gqONtYOzNy/MePY7PUbk7Db
nMJXzMxulQjdH94yvd/CyGHziEvTTTRodlsPTlJbIfh7R9gQTujX8syb5ch+Bg4R
bxNACWtFfsoo98Mqp+cpa04LN6M40pvuu1NX3dnfxgQYTVfpLsdv0m2wtlpiRBIN
cqKaaIT6WFg69FRjj6wATWcvqBeRCovZQAJBqXNTkxv/kCof8GPJP5lysyBU+vlR
sjhovKpV2SCE+LRYcK3QXJzZh7FAuSFPHEUzXHrSsfnw3Q7++8DM4I3XyU1o/lLk
aJ4ciaJNATcgil1yjzL5yeIEnH6vRpdsU20zrNTaaQryqOW0lc/IYJcuVL81D0IX
H0l/wCJQs3kwtqAEIDperAo5bj0a31K3k76k3gLyyGMInUYprI0UjCRLoTCRpXI+
P5mfPj0oF+UZAJSG5crSo2skg2S5mPIzX2kypGZ/ey25D5dsbEWD5eF3lswdEfF6
1prDW7ASh1buScNCyrnqbvvxRqgLfwM+Il372MwpsWtL65qGvc4UwvUCJWFYVlBL
JVGdo/ABavDVWM2+Gkm/vAkXT+i6yCNxfsi4WzbhRFXM07KEGnDG25aQH+0xW8bG
U1Q59ok1dmVUwV5L0QBMWBMp74m7N2juZkV0Y2qe249aWVRGydsjJmc8wJ7ou1Ls
2JldTAvq0u7pCgjA4071s4uo1xp9XzIIimwECoz0Qh5aL9F1UYpa1+txQatq8yO1
ntdTkXIljkhivhrOME5w+efaTlCGTb8CMG9mNQc+kDghwRJTEqpM/RWW/lQ7Zu/T
xboanJW/44t3I/ah0fFRGFG2tpa1/d38n0hfvU5Dw0K5LYfqP2tpqNd0Vn9hUsL4
vo+7y0TmxEEVwcXq2INfze5YZJaW/McEMIOfCVrl6novhIGTe1pzr6tJX2+nw55K
quQCnKU8huclo0CnbqZTXe3pLoLDmZsD6BjtSW+6QE0FtcCEJ6bz+4yLnM8k88bA
SmCri3w52CRBoljQM//Oh2kNEexgmWXmAlSD5RJKiAJIaQOgo5unYU0kYfZNS9Kq
TryRVLtT+9cxEzRDaXUjd+R+Azm1sovaYsPVZlr+n3am4oRjIjIzq6Ng3smsh0bF
FQDQfETFX23p8fstH/fHRNjwz0O689dDv20sJsQYlvRb2JhAVm3o9YsQhvf0KwQs
JDjg7j617PBo1HcdH05117zHS1q/9soPmwBFL8136WLHzWcg59DTCa8igjBZek+r
WoU6nsHsPWG5CpxqflpKUFAK5Y8MZAu6rxx18Q8/CjNCo+L0mxFfihCDpkSjGCLH
FkA5RZgOVX4zBQ3q3lhqSoAmyWZhzB7yyfMV8Sc0uLUY4ZiDt20iOyPLoO26/Qx7
y5nCRFZFVRUliXVMW2RIygIFSHF2QBokpwXFFhGn2CcxUW/jms4ABA1GUxv1B9BP
ykJRRwO9PKX5wwRkqY7+wCxcf9DsVAMi2Tuv2guLTwt9ZlFzRRHNF+8ZsDtEkMNL
yBae35kPhw2P0Qxh8n2j6ycnTD6xJVFKiW3dxgMFGolP93nvHDz75++e14Wrfxa3
eHpOGVWKjYWtNne0Bu6APDBGopzG9PRXIQKs/HYPOyeAH/BD1n7kjFrUYPP65mTC
4yuM4h6ODhutAJhfUJ/QR6MRS+qrnRJPLCV/Byc+v3474P2Vn5fVmSzJ46QIlB3C
K5w3+Y/SLl1AZhnrZgm4SS1FAnTXcH4t9p3PHJavYfOyplDHshOvT7116DfKXXJT
QBSK1Kvr5bkarkM5I8DGQeSp8YeniMPACk3aKve96Fq08zHSGW8ChMZExF4S+OHV
PJafoYEKeN/p+qRAjnysdsdTGBXguTzevIoZofZXTNggEax3IJTtdy3bAEQOz7cl
djYoK6138GkX09En5gf81V3Bw8PK1+/aaCtbtQ6itOEDXSKhiYKtR9VxkLiuQsS6
R0rgVsKR7a78OkQW7Hs/zhF3t8CVjbnqJFUHfqwErHugyR++5X5UiE1WWLSvs1cY
9QLQUPgsE4UBIvysKPue6qE2ooJJFsw7ALtxdNjE0rHOD2+R3g4SajO/28PteWPh
/2TNNZJL8BcVGUXDcQMXRL51DJXk/fBKc2at6ZhXK++jg6nMJ5MmPNbyZN/2t+F1
LmxTL/2yCKeQueKC/ZPSq7bveWipgJ3dR7LJ92ltzI0CvjEqzfMrv9mjrTbtRHbU
o+wLiGYp5yPbdvG5w7gDaVbBzc4T4vEbpBdIgdOqehysmJfAKeyGpQ3LhN/afbGL
yvzIFrhpeCZU4H1jMfGaF1h6hQ3bjIthAxpmWb1hojjDTFMVgJBwt3RG38DLC/Fs
lc3lRXpke9FrFCZWfFQKcyN2cupalcDcS948Xe9p2M4vy/T3JwHIgLYdJjNfGxQI
vFHpVdwZwvz0YRCR5PadcADoGmZx/BN3vVIdc+Bsk4I0BkN27uGpt78bc8eg5iJJ
X7D8QUVG5y87JNK6pfkTv7XoUhhXE8EG7fdX7TjER6D4zW0QJR00jFQtsQ5euHjI
5L/X64bgci+mvykQdzU8Ji1n1qG1uoes/rOIh8BjuFzveuBnsrURXFA4b4mlA38/
wXmxuqwpLpiscugwINTeTnXSGHwu9oQ1geqI1EoVOFESAxvBH+W1l1UbAMTCOGQc
Vv68hduAI9g4VScR3MIDo5e4FS0qf//qni0AZGrGhhGzITZs3FUVEIKQTHt6QUAj
mcoLlp6B6a2JbdS8kqJywLlzS6jROAGvjU8oVTE8UtJnAooHIsZ59Ijkf6KJyN4W
nUzzeguMxqpXPzBoMPP1unPDbEtvxT9a6ZowOufdgm+55yjI6dLb98A6z9+Tw6+8
K9Baf5X/D6eHVu/jdNQuTawZfTL1H64B3LgKfNeiw1520nIld/3F+fzLKuTX1av1
aAQqKmATmJcC3yz6xYhU1HiN8DBqUcqWrxV4nM8uhFIizAgpZniEd7NeFh89vzjS
CmUtg1w+85rfkfxRv8GEG1H/n51MisG/BVTUjjJ5Rz/ksuBsbqEF85U9VPbn5lAT
rRMwHucxvnw+HhAYw4fNB+v74PRT6mz8TWKws2bf8lIAMi4+36FJYoEJt5mGsh+p
cYDbRvYxXb2iTXWduPVkuz/1k0V3LUUxaYryKZajVhH1UlcMAq76VPa5TViGpSHd
PxIT4xm5VV1rHoRnfZO5va4ueTlcmpWr8rdjMdFKaBWz15VrbBac+1EHGaHV3ehH
kQgc96Xhbeff/syG9/xOYpUteYE1OsDPf/miKDoFBifD8xKskcp31MXNIAlt94KL
WU6jErqIjMJ0AM7lwBYoa1E3dUs2JWy2vQOcNP/dGwM8YR0HWnUjitJV7Hh1mevk
Jrlz8XVhvJ0ESQp2uUXbDfOyvqw6StW3OIr1iQnv99x58lZL3RaOlR5Pa9nVKeC+
Iq5aMv3OmpGvgnA+roNHPQ03dDBUjXRptkJP2Ozrao5cYatF3/cQId3v0yG0sOtc
4reB1tF5a3ILXH8hK/l7J6bPsF0HDJZx+bsgduL26r6/vlFL+YQODH8yucGOOboH
TeSLEH/q9lkHRL7Agkyj/kn9MifHtdHVAJqNZhsimS693OJAlckY71jELWfpOANH
Ufd/TNRGJ3rXVZEfPNi/nA6CvJs69crMTND4ClAsDJPcXaQLSDlA4K+Q5VQtZrm1
hPsEs9b5E4JwbOs5QeMLK+tBI5icGYrIxzonWEnUV4jHGebQ8o7anURz0xIotUgL
LtZl0gqc9GLgG9XQCweTap05UWiuDX1fMJkrsgb4xbvE+nFfkXIkRqE74GpD/X0d
s/gs78zjloEycVyUXEDIif6uG1tLvVWBBDjFds+8QxoEDwTcN9nuXfVdnF0sTysU
ncdYxgRts/wwTFAWJs7w3LymE5oy8Dgvsj+/sQQ6lWodq4EMcdKyR/VilIfGhxYh
5KQk7982MOWwQ1ap/rvxscHjxXSMzjYHdNGBYPnVnrh5K4IkwSnjn1fFiqFsxgfB
jnRdwRioZSndPMZ3T8/WjcgDR0OKhNrV5+6cJf8e5yMbTutTda3hrUzoojR+2uBU
Wp+k0BF1iCK+TTGM/0ekf8Akd5nVpgr7gTdGt17IPjwXHsYUj/F7cQ/we54nYYwi
iEOJI8gyeP1YcYwiAHcDWdfhuhgxaXxw+wkK2hX2iOIRuny90YSScaIqKj+tySpX
2yBFWdjzrQNaS5tySx2rEdon2Ub6dklPGfdU9FTUkKkKtpwNj6fP1mFzu9TRNKou
3m4Alhrsbxj8kFhAPGFj2lKc/eoisBBOrSgutRxvzVTdsXr6l9WKOb22xPyxwaNY
uRNxPGcGBkkxa+2kS9mhN9ALqAEHA2pOxrYAW2+J75MYzDBE+oqhSoiPHxtVHQcU
HLtmtPEsoQBuWhSOWhGl7XgJcMosUn1ypTikYlS2CqRQT7BVxvFY5xtUVizkyP1X
o3M2o4Wi+1UMgpQ6E/ELDlrwGY13NEryoMFGDJOBC3mlE/t9QhxRrZLl47yhuB14
2+hpiY15Orfc/MGCafaaDf7MD/BkotCrHDULOWskY/cW+Tq2/IyS1jHdXjluGR5s
WJNH1kYT7qql6xlweq9p6WR9vR/F6Mf0FMpBo6FvPzNq0Csu9JX++JTDjqB+6IHZ
JfdHGXSNECIpR0UxVe4Luc+/TMecI0QEfitIpjGh7E9FDY/zAAbLXvwAFQh2rd+d
Wj8RNLwAnKd2nKT4NvDN05+pfxXAYsADmWSQiHvTHXVGYQEaq+tFH54kEWTWQhGz
u4XN2h6g9dZekrePML3xX8/zyJIdhfXEac4BIzKKEbijCPkoIf/4QnG0qY/KNLbf
jgCza3J5axmqdcTt/sG0Os6M38mcfpudU/ERdNh+iEFHKZxBb7oHGhZrBrlFQxQY
RFC6Nck+X+JahMsMt4iQZaHc/Sfr8sPEOlqOBjvdELl82VoA658Bk8zhnWlKP1oh
k6XQH4IoKkT1sfhs70UxPke8yGcmkE5xhb+xi6NtqDPfxhIE6IGq05xdXJXrfH3S
nB7nX0yGDcFivRifjXGgVD4DcK5PBEiKVlKP142BUdthbbtFJ2ug3EDQcTo6Zzb8
uRjLuf/eK1l2FkbIPSf2L+ACN7GDnLLM15lnBaaoiUBgvcS3+RO3p57BsiNDvknP
krga4UgdivPxlrpXxs+dHexGQE/IhMQWKcUIDXaIIeHMh3p3xr0rSW/Y+HOCL8+L
KfYVGnS4LFq2UopFXwWTYLsmCIeBCrVJTBPSiZl25C+xQLZNNyeMK2DFx0nOFVUB
MAJCJuMOQX7Q2OShSM8Gmn6PZf+bZOrIXeDld/Fgbcvfr2cVDV1/yFwX6ii9EzP6
OKou/pVWG9Kys9vhZNtTvsM9qss8RoChrKZ+L1BQENPHn/kK3sJcZtUKARtKsosU
u3p/5rutVWmyVLa/3Byn2dEIguQimZ5caoxeR5qjYlGIPD31WtRZzZzga/w2yHBS
CnW5mSTyTxugdVdU724TmJTvcfk0n9KwODFYHdjmAqCQz7zg79B3Rbo/v5cB2dpQ
TcA7uhA2HXlo2wwuCVGG18MRgJ+EUHpnnCIsdvMM+9Lb3BDaXHfMNPJZ/6SUpVv/
a8mWuw3u6l1p51yw67YoOC+cRtcdIQy7O4SR7gKyxf6CcidNdRqz4bT7ZxL88wv7
n8A8ZaoxSRJ5iavQXbNuh6wHsdBuYtSQecXUCj8jSD1DGkofr1bey5vVnaESN4F8
4nr6gPSDudFB9acNOPGU0Ldl7u1Q0Dl6Mm6F4blHOE5kgFoPo5xS412+SoChFBi6
Xdoo6ZrqXzgSKRD0j5F53iKksbm7hrQ4tcF26gYEPxS+9I3ua03K4DsclP3VZgsX
pOgkhGcva0vNFQh6Og7YoAgdshZc85y78iQCy2mCWJtSEUo7+xsDks53siBz/VKW
w0Nxkn7Tmp5vLOZDAXZwXzDUyTCquKW93YK7t+vMwf/4pGqV+Ij+3qgR74iX7eZC
hkcVuFKet5B/0si2dC1kF5kxjgx/PKLDXHjRpyXI4S+L0yxEUWxj/b5wngtF2TJM
groN/CrK5nM9OAnsAKFSj5aFxV00tTm7FlMhCh9gjBH8h4HcpTNhbaenm0DISUtP
pDfnIB1Bkl8RPWSCW3eYEMTbmITPcTgvL67gPBsOH2mcWk+Ew0itedjZaFzswXSy
lbxtusgZ1GfSGlFf1RdNQtV6VlP6w7QG36JJE38NhatZt6r/VTXH1dHxijrkJYp/
LEyUDe/0nIHUDASzYN5Y0brzeOu8eMqJcXfx44r2w4V0/sRYi2p9i3P9Iw/UfuzW
qzNZVeXzLPvn7kZ9CmonNLl4s48kTvjP/ZLb4ej/flx0t7umCs4UJNWclapfu3uS
ZqPdbUQihsf/dUfw6wDmgy+ONQrvSndWcP/DOTJyDV7nZORwnGTi/KF4wBQZyCbI
4pIKYZzLzVH5HDjGgRJ1kZfOZ4rlL8fw7jh2xyDDSKDXiypNvHGxCyPchxoq2ZDl
Ivdsr+Js5orT5PW+YC+mlUyBtJFCMD9oLzpeoqZzAHOU9PLBzBFanHylirVNskIr
FaLTLN1TYnJcnRLmph+/ON6/DcQ3fwSmRxGmKPq/P6aXVp4iRJtZiF5a8f36Mz1i
Ke29REpK/jz7MbQkFBd5hiChQsmLd15ujebUwRcI4TXM/yNiVUgEmN/hWi2kEfZk
lYu5a5ZxJOr/DK+wOFWzePWHDxpm2VQ/k2icC5EqALPTbBU9zBgzCy/HIM9ia0CR
R6HZh50GOEzaxlMC5Ha5uQDlwLXQfjN8Ry4RQWmWvZ5qvj/wxc6pG9uha9mZsBxi
1Ez4EB9e5Rz5X/vJXEf1kng6ByVaJOft2zqVT5lJ6zEOcfXqR7S3CzBuRKV2QluU
2HLyswguFFsxpg1IZeOrMSrG2ZCs7fXC/Y2C6O2tO2nSs+VfZk3InAou5yT2czA2
wmWjYbEFJZHhhdpaVZ6cw/oxjOk92VLjTtg7z6Kr/KDlPl3CXPM+DiHxmJif+SNS
eOekAsC7eDda+7wuqtF2dBmz9u5z7b1tELD+hIgQwgYAhxP1V4Hg1GReM2E8ZpCO
/z5BirDkN3duLtXUZ7qv1k/y2tVULhjdpxO5BIrNyR0R/gOU8+dwrArMs8Pqi7/k
+NI4F2wxIi2O4J6Xptq73OqR0UEkbb0jpJ7+nnjeRUfZ3c3lCqPFwwfRINL/4A+e
NIe1/SIeptZfzGsBKKbeNj2FXUEolN53sGvvs83Xc+lSuR+gvn3k1t55+ZhZ0Nr4
9PQ8XnkmhZwYOgq4XOx28QglacUJYUsTm6b/Z8dvw+TUauR58SAWyxApRlyZQQbo
AFocldYFdw0fHv5HgVrRqubx00XfiiKR7YjByq7BmuRdFwgUWCCrPGO1HwVbw8WZ
B18YOBCqie6AfIIpAQLKbSBdrSk7Lmyq59z8oFfJ9rQ/BwMBsrVBTNKXyXZprrwv
/gBp+cwijYDxLHKbhOBRpUlewdDn6MXv9J/c/E48IIkOgsXNvsSKV8CFk90p2VaI
veuUWxqHeyzMasWkElZnfr/jDx0F0909tuokQER7tooSAhqZ68ikW9FcTEQ+Z+ey
DBseprL3riKaZ04EAxOWuGr13yk4G6U3rjrD+IPKnH9pN02rhMXBLDJYlVQjoQzQ
VlE6EgUAEYVF/xpYSU3lalSXoiv6HUeT7n75zt0GHwO8qDUCwEJUES1jPdvZ4HW0
J8mbgB8j95gIVUai7sUgOsZN+hHLhpZQ9DEQeQ7X3d0BWCSrf65QsjOVXBpuwA94
HpwQ5CczKtETp5LLoZ/68Wt7WmeiBSoJG1z1udML8D1Ld9CsnZL2JEcNzpRjzjmP
KJgSmPbMyg582o1+r+dUdsQipUYlvgvBbQ10oqJGkpbT/JxTUS8gNGh/2Muh6lKu
Ae2PXEkYE0Yr12YeTITNKZk3jEqUvl8Er0fSJuii7S3xGHFI8fpB4rGiJ1qtnCvP
+t1eBPYD47E5MEqsNxqLB8Ig04P4ESjBamF3UGg+7lACtgXTtRL4MR2dkJUF40rA
Yxu1gjGIDvxpxrK6IxMni3UZ6OLEYktY8Tn0ZcG1Cn37vfNEaR+vsb3CNOmk1iNi
FJJGZ02tZOPZOMD5AKNW+Y4Ad2CDhVBPsaeIgoQJq2M7lGrhqUecMNeKJZhXQT/j
d+6PjghdhBVwSHK+e6Q0miOLJSNL/kgNWVxkqaj+1LXUqr/+LtPaLqxVkcwXq0nu
+nxF0bqjfKqS+k4oN2UJ05xOWkicFEKqnDJ+c0Um8i8cMFyzqWgrgV0riD73Dxb9
X8h+rxvoE1mL6eJG5TkG7LmGbGrM7e4/vCNIks1pYSQMlHFwf36MsON94JM2NZNa
GVI0gdXXKimns+eA0fl0m9ROxdr0HfOxUS3KRECzN/t1fVy1ABOwty6hjeElyOPi
J84KYvdZjWcD5/QusS1kP2qwefIkRNNoZYHPztbhWg2Vpi+IyotCW5fWDKubggSO
AUNLOecDRM+4Qpsiz7+M5X/9ty4vxJHf8uq4Tkta8J6S8agMf4N38mxZ/UCZXcwY
Aafe3xKr4ixNGfTOaVcaUqJDsgUOA8HImpOKFchhDG0ILy2ajQJ+8DI6uC6hdsva
5Vp0DwMqqXS7zGZgvlfeTgR77rvot5AZWPXhGf9FssJ1ZM1Oc5I2/jFTEHO6yd1K
LLKmDivR+/meZu7+w8RLUxNuJ4gVnMxRLYsTBnR2Ekll4uvm8k1qSNDggLx1IAKp
4jNb7Dgw3mFIv62GqDJ8JcOubh41j1+cadFUFOlSsTIMimTpt7XgypqcsD5ZdR/0
N0ZC62ntpSX7HyGOhqz4pT+ri693SU9RpphgaV+yDB3IvY0r3vOciQozJfy1cpo3
/MrOUTI2vcNzJeGWHUYt3dWb/GHTrKvzwpdIIW4V6JnHHB4NXHgmnuSsKYkt2yNB
IDGmm9GU/2rss0yFdL8vq/rwFeuh5TN7VBcRtgWQ9e+LhLmQlt7wzvYEybWpEJwz
ywt39DWPqVeO9La56uaQzTDEpUhjq5oEKUf+c8092Tr8IOm7Unlve/Vx3U8wxuD4
csg/rBANdirDVACoHy7PcKYvM6TFw1QZzLeo/atBP+KxaEn16jV3FGY4Tq4OOa6l
3FoirZb5ASh6ZkjAj/BqgeI27OXWhM0RmSQcOemWMZy1rWQRzwwedMyZ0sLVeIZS
f8n/cqzEKzOo6rsq2elgyMyspesxeGbVcdCouBJl5nCCV3+CWTkp2/pOeWnzEFUv
o8QkY7efIjV6J94rJ6nPfsq7IfEJQkq44NpkZn/FKIN7FwYCcwKwSiA4ALU11j2f
aXpf+KnAbQZbRd/Q5WDg1F42JyPJioiWLaj/7jR48EJ7oZE4X5SKmrOpyw2bDojE
BOQQ4QsiHg0H2A0gFTTFCPkFaKcpOli1eq2fZlk85i/vw9ryLUKtsnvvgWDhTuZI
fBQBVutVh/RJxx8dM9NlR0tUgxiVTAFMJOBtXydX4WF5tYRTqI4uaTTqpvxE3Uov
muPoUCSTL2h6CBJZVsQmamSZFhgPfYczdAc124cDzPOHbO+VUNp525C4kbML4Wp2
MFxxQ7NoH+6t8EvPANyvFwERveEYI44ICdpS9QT+jtT1mJmMs3LvWD262AGmkeBV
RuKmyX4jYc2bjXnF9FBJ2APd8MgxpydYcX6ajIyuBT5n24+RYHnhufkjJpWKpi4P
+FloyTCozODyWcH/qndM4baKGUBZtX0HuF4VOSafqVActkH4w6781B+C0ny6ua95
ZePrdDUdLWnocRTOe6CxL+cKII2OYqE10pHudUxMokTYj+1zt8B9ovGkRntxzWp4
P61uI5A9OPeRs+eG3xz9dhoSLmjaX+8uhWCq1bBhE+10lNLDoVGp8Y/ixCeo37qH
tjHkbizfpoC0ZCh7sqR+1cG2Wr0I4o8r/wRWdYi1KVE7Fznj+eg7QDRjEmHOAhsz
nNJZWkPjI2b+ZVvxzffuDWUnnObOWjA68+Pn2dS7qk5PXVFP68NTyXIc5gqT2B61
ENOCBSCUJvm+3B87+uJurtjLE8LgQgBE8II4RfXSyjKW8V5TEFXrAMaOCQFpwqET
MozCftHEXQguaZDXU8JX9NvSAlFY9/SoD9KeAG4gsgDEf34UBzZoWJWnXu+PTjyJ
c7cl8W0RpnLls2DskgTRmVXdJgeWG5ZRTgqkPapRQEwP5QerFYSP5NNFxRf78V1Z
PZGh+uXvvRvqwnw3qDUZQH6xoPi0zOzgjqiREaK4NWBRZfNq5j3vhku3EgJ0E9ar
faShLyrz1E24iDN8GsGVZaCIqUOiJv+sTyd6BJ5C4Ap0F8LTczIGGQiX9PnDe25d
IcgqYzk+ni/kuPrB5aPJ748hE0X1YvwZQ/E82h2CRK9VHgu9eVU985dDviig8B8B
XJ5XlRG/GlPFsT9on/sgdSv3nDqxhpmteh8RqpXlP37ZKFx0s8H9+oJzzeLLnvcs
rH/AeTR4mIowk+ax+Sz2jbKqTLKJQHzefPdkGKoCZH8dKluplqt8byS1cVWNgb3M
skleUWgdHhQKYrsRO+iA1uWtfsCTEOlOjCKUskjBMU44tLsh1YMsgTEjOtL+zSc7
UTVAgu2oWTypcMc9Iz10uArh/sRnLhv17XTq7ymycSxp2YEnz0Cr3PayQsbxQTBo
MDdW2QAwjQZkv44krSJlBZ0zADHHTV9a8Inl4rtCTqUQdo36yrnTh5jEewFZQkto
kf7YN5LKcA6FLSBjqAaEqS0gdKbIrE6Ok1SEgFvdRGtptPCPriwATMRPcZn41/WA
U0vKghJuU3TVt+4hUc3s8WuOTeC8Qg7nigVbzHg6eVDRA26tLF7Jfe275+jBrVvQ
vfNt2W+uc5NHfIWiWp8aUPTpgrNIK1v3oTC2ied/ky0BJqxziAOcLXGoQsSxsrTp
9pqu7F7UKPfp4WLealVeEorHAOIQnBXK4ymGfZACC6DfSm8UMpSiQseOikyeI40k
+1S1e3jPo7kco85u5WysOb2gIJQhrwz8bxeXsP4loMsk5eDW3nzTg8UJ73q4taes
dIGpX5zkk67t1YSqExdQURbR1bxWDuyebMtpAEPNcno5ScAGKcJ/150ho8f3zmn5
77EY9tJfVYt5zrrVfbAdfEXUTtQkUMLmgGaA08aXIJFAPtvhYjrYtaLZ/SBJL9xb
t9CsopMVqKDdj9/8EZmfKEzYE8x/67S+qwAcB4nBLHYf5ZiABi3wrUKQXybxgQ9/
0cq6Z0g1klGSSb+XlA8Kfns1s52VmRKsn1KrVCnUDA0nK1EdbviQh9erbeHjPIwX
VXr5v1hIJtCSMAIyNphc6X6RldrJgFqKaz+YF01Apdp4b+3JAW+cqToycQ/i2aXP
CNFEu8xhSy+Uo5kXj0oCL9dBCD0RI8BdZDIsRi8rUO9n2wI/iS90uE4EJZf3X/H7
BKAQ9EFUTrix43rzPXA74LjOu17yBhoYDI4Fpv6pgGOn3rnzgwch0issGRCD/EbL
j25xWIMuuvZ5Ogm8eiQMsL0mBZC4bQ2F7ty+LhaLIC1/hRf41B06nkaQtXY68yh7
28qzIZxUeWQW3SHmRBi1RGWKOcW2rF7+MFYWLrdlcgAeY/2RRJ5KqJz/zRhSPJiG
EQ++eA6wiBvMwYIS5lFWa2zqy3ut+ST1uGwx2ITFLn9qnE91yksgObWgMBr+gBao
xRTJDww9jMXL7CjZwBhQ0bMe1pQ+iVNIOhgVyDfoT9LmZcnH+9tJOaC/tYVPVIgo
4/Tk6mZ17eK09KhrxZmS7yA/wfWcR6x2UbISo1UBPgFtMA2de/OdRBT64FBn21Bp
6QOCqfXHZvFFBWJrhN7cSaYQuNOFdsqU957zodKZeSee6EnNOq51T2jd91xh+WmF
skjcaRisfxsutjDKaLE+yznsGaLlF8C1nhy943AygV5wvO6YC63SCGp6ZJiQmZIY
aFC6zah9xPcg16BZsEHsaBWlOKSwTiQLfqQfYCiyLm5sgkU1qOL7hVuj4e9Q038p
OGoRhgudI+FfrLwAIiENMIUQXU+n8hBQA+kghagwwm9v+hvieS3Bbc52HaCury+7
h6AUMNf5Y/DjAFCtnKdLNxVnqKn2RWqRAT+boEfmOVI0mVa+ZiEHUFRg29dIv0dc
clYDt4/tdJ4HJ6toV56rvfu+nVkmjWKaBbuR0HYqB9m6i2uCPfgnh7tf9EB508nm
+BASs2z5XccqrgWGo6qHvhhL4BcL+y7x1yn1VIPdCzm7iAtB6WsRR3vc7W/HEq40
DMKpNHub2+WHrvhjAjW0RX9HupGFKmM4FwiifFQgPV2rY44Oz75jiRup/dtm4npi
rpPz6XoPXmSYj0pghy3hZXDYPCCGeDd+2P8p4SnpBeW54q9jJ/P0dOa/4hOeLYMI
kAHRcUK8CjfQKj+HqC5zAOLyxOPP8AquKj6Uj/iJ+uDUiSzxCwec0wXugZGUxIRW
ZDDQTSBiU/NGkUP+6p/l+Cmwm3By+pAQgYMgXUV59loyPvwH2n+zme/2Vap89JLo
T+aWnywOa63CjJU2fFe6eraHTrZG5VF5PvXyumm8fbaPQ1MUkNO9cu6HQAXDFO0J
f/OTaB3kGVHzutNnCU0Oc7JhMB1F8jxEajCvsk7s0DcWYGPEpPEjrp9E1+chHuyv
xl6prt5p8HcNOeGDHXo9bTV8lKx/EAyC8/SMFrU7y4kgTPcGVRTjFSv1JKtrtwrg
A3hf5RpJ5uVSsOcjfwryvnjuMQhYFR73yOtCKRaBmviyJVvxoskqkR3ZOpTSMjZI
06wcAHPBpZl2SEXuNN7I6Az8LhGYnVnVPPHGfzeavEk1NJ+Pqv4EEh1OnMAaWFlw
/3lr+8ZxMcoFy1QLtCrl5vlapWwyagzz6cWDzvfkFDwt+2vVbKDHkcLoBNPSWRgB
eSroPbDUvrUeD6kc/AfIr48y/AWBAOzUxI6+iFY593HRDdavH2a5LOb1VRWU9Bee
mm0NO0grVJGJoXI43t3D3vBkW6faDHsKMJL/kIxduLBqnX/emsXRfaXrwF6O+67y
vN9zfGUZA11ke+XrRsrJNVMWsmF4EzE833NwMUWDxetI8OLn5ZZ+lBJQZmoraBBY
/AvZqvv/ZqL86vsPBE5TkyIAtmZFu+ien0jSwmnjSrw+wxQ3cZDyH9YZrAwgvT2Z
H2WBXoAbuwXkveOm2VMPNis8NLTDR6r3mX5KTOD9Yo5+gOQEQV97VsrrNBV4HSXZ
4XDGc72N0AeSRtPK0VZy5NtnbuabpywnoD/TqUMw8ZNyU22eCGJDhyTsifSfIpfX
Tz2Dk/xTEOFaYmRHkYCTWDzL/pK0IEr4JEyo0B7xdk3egESULoZ5nBH+Ul2dk0Ow
3AiAE5vjsUNiJmr9fCxBLdBBfhSfT8WJi1C/ZtKSIzvQO/C0D2sbNxJvNy114YN/
Ka8KJ5/LU5PztLpW8ZYxWNZcmkUM1sC8Q2y8FowIF4GbZ2FLe1STKb2qB361Z7Ki
i1tDO1V8JEvyFpdArQNavixLiEJOvihUVZth1zxii7iQZSSDv8Z+hsH4xWkywh+z
lBaou/6jCxxaQ5QX9rdzvAFHHLc8tXSQfaWAcYVYEm0TckbELLhhRjPYqyXfJzuS
oLNg8DBBQj7Q66Q3ilEeIsNhykbsvTQZrsh67JAwbuy/rqhtR6T52ePalJ15knks
BGR7fHSO23ZgTJ/K9DugBmfL/Xk61scOIZorK9ZyH99SyfzKpL7aYMk3D4xEzZb4
k74u2LsCA3lhzDz5257WgpGpHnroIeK/F4eFn4imv8xaoqnwle722QJfFzUuqrRV
gswPePrvvzRA+eFFaTctttXRdkddodV4NLQCeeVa5GfWINdGHmVOr7E0ndn57KWl
5RUvEklA8qGpwc8jyP0+/FtBdPCl9v5UaJwC0aS1Iz5J5IAAt7eY2IacYA/JrAzM
qSS2vMM1o4xmRAXAJNZbtbKa8HDF0CjdHRcWfozjhnumUDV0f1prU3bn/81vEnY8
6vcgOi597PVqv65HMslfZ9VYLGxoH1bEYhEIJ43XSgGufJAdtN0qu8sTsiFLH/Su
lyDZ0uRav00cNEojmbvB8gSkYYmksLPTugQUgrDvCC9xD6DuxSbSCiuxAAGhgfqK
pnsaViOd1S43VKc9P49SMTlzFnD3GSn7OaTuXGc3Kk8kmGvWaGPrTsnSxVYaFkoY
GlyR9n/oFr1FJPSzP1mWQ103qatMxyv1YZ1OlfoY0v8YarUFJRJO9c2LCaBBcgw/
/jyrwH15hptwZuUNBWGwVnUTDU+K8ay/VBCCbK1FLo4OFg82GoYSDHTXeLl02Lql
Tq9YOUkSAYjBCPd435jBApUvz5zB5zPhrppTZB6OHaSAh3OJltQ4p6J7w54eF5DS
e5h3RSvOOtG2VK8AxzLFy/V9EXTAq3Q/YEws2uYaaXhAlAdcWbML5rzyWDlY30oF
forCrEcYITTBpv/UvT/tJ8s3AUZYUGlchMqP+4yEbKcb+ibn404KcZ6bbD5XEYsD
Vx8wkdoQkf+Ok/XlaO9Q+kKDsTTDNVqzZFommEm1BXXRdJWr9sgXLv6l9evZMNps
uM9oL7m0MXPbpgpoqiRC2GQV7wntlOIud7RY0fJhpZfQ4UUqo7h2RWDUHUZIF2hw
QibMHPaKCN0Ot/1jjfwqtv9BC/mih6hdG/aJEGhY6G8OQFVnUJuOtKZEzR4vz4gG
HPyVfCnFTJ2dRVOxhrBT+YHYsYnPoCk2ZHPCa58D2x4VJVtkkNvnsCBf96cr8p0C
SZTCBDgpq0QoRcGtD2ksutKYuVHOO0MmpLI/l9hBAu0CVGqaIh7eAgdFWybawGFX
/ItByk120OHU9rrqXtSFC4XEF7p+gDjzBF4hHid0mcBaG0DZ3ND39QFRV5jfYnHk
JPxCYckRzord5TAhuroFYHF6tNEvZW1hfgQeM6tk/N6SWO5IHmfODsTZe+K+XtaL
/nvsQMntK+FB0xR6C+gsifPbJA2tczheAx1TKpg4offMR0A4oP4PIlYOyxR1ojNs
ks9E9ivcJhk8P7Zq47Kg6wF41MVBC/CMrRt5DTNIoh5agsX2AUOq3qLq9h6SvicN
jT2EuPCVPEwQDglzgUzSZYeqrzFU2XQkaHwB4d2aVebKcSoytHEJE+nutlqmTWzM
lOXJeD683plCMzy3wBjF/XTGgaKgZYjfqee2L2mwGu7FWYTP9Y6H5g+WlI4gj0od
/2EELInPJXibbSrfM/NW76JdjjnCXHAkWtVAKQenTEbKU/7n542kOHzYZmkyanXD
VlL/R2fH1YpYagJBzfBafKg7yEYE3tE1Uq30OsYGT2V6C5eqzoG0rD9VFMvcYvWk
kUp89k4Ba2IatsB3fVW8/+SBC7X565QJMMFABBw1prgJFYmaZ4KPek25G7zHgI9T
phRNw55l34qiPxdTqpdbr2l6+BziiLdFFLNFzCr1+XwfNosbiWrSU7tCoSTCkgGi
gkYW4FhlGq9ciOjcfufZlBiX4vd5L1MYKbO0Fr4pKexGQcRvpmg59CSptY9b0j6j
+JZmYAdzKF5pv5l4y7smhvYUm1T7Mpla3DhNvi5qahVrWmO6dKrlf+E/Ybm2THqS
xsskAb7eYdiIRG7jx5FdPfluU0xSW7+bCKG0hUAi7Wzpj3rmUtGYFKP5PX7PFrei
IoWbIPiuC5rKNeNceAgX+FxTv/zKvF9CmuqfMAFouCE/J9wa4Qxq5i7TG8kaJgmg
qmMRQ+KBG4pXM8VzLdID3bTY7qw3XgR7H7oSTfaop8fSFhf6LxXRa3gkbbjXwFae
ROIiO8IeBVZ88AbeZFE1gRAbez/lsVy+AepPhK3TyORVutaJ4fzrN3DFqORC//dR
vreaMdl1LstMUuGa5d2RMGaZtnoaLzQUCLGbGDI5EwfivCCbD2BYAGG1cVP/zvbt
mOxKK/vkeSfqGF/xHn4QbBUpW6JpmIiTJfNhWuJN2dfP7TD9j6HgH6aRcSrLqXuK
wsZnTal4Bo5irs8w1ICmXZOfNNpnZ2V90T0Bt/ZhbYcn2O5Mpe65aXbMWY60qCJK
qJuJcIOi6g1m+pCOrnlya9G8wOZ0v5x0CxeYVcy0lv+ckvcWXoXyCI49UoRVev+V
AqLQkD/vWimYTuV2ysH2XpBNxVVAyYyu0GS8cEgu8djf59xiiKbD125MKK/yhdSk
HC93fJ+jSodPIDREbM2D16Z8pVtLx7zyF0KKTdSIB57XkDiPy9aTet8+5SC+3kuo
+UBSLthhcTmrPdEWWnhnkmJQ2XPueCSiPsB2WNYVH4onU0hktgitFzNM767VAbt1
QFNkgagrSmj/UB6tSXk7FrANVqvijGYOv5mKmv3k8AToLo8q/rqUGqHW8a/gF9mU
Bv9MW7OROETxRaV1cne+VGJlpELFqMNrWGoSKT8NueN4IF91+wE3uq/Bo65QroSQ
X0dlLxKIzvuqGFY+QN+P5tDOm8wfaduMU2sXtISVBvYPEo64oyn5OxM8ao7rCgV6
+aIYyPC0cBDeGsqSHeg4Oslb03eQ6HpUO6N/x5hON55GBMxehxrm6tkqz6BGZRqt
oP7nASkTLu/KOIYPbEjmLTH9vxY4SlzhbCnP4RhJeGgpy4Tohzd6gbAUiopuFoHe
3z7MH9lPDDLWS54ElRz7Q5wyjlihSilxCW21OUGn81z+FuU0XhTWN+cX5yeX/LaK
nqQDH+DzBgA6yhR8WkAL9kMWbPmtrFDxdOlP0uPlZu1iSVYGN3/qc1Qd0ILWlxuo
D7FjBguHPvcraOxcerGK/dOZORGM1L6fTqutg4T4jTNX+ClujhoQs6P/51LeDrzr
wNiRKTj8X3/oxV7xvHv0UN/U2o+VXu0Xo1SaVphmtPfC1hll+CYsWgO0Jo2S16g6
gD4J5C4HmdMAmE2Dhf4YIyOvJUnQHeKk+do6d2eJLrsxOhp9bGqhuKj8b9iCuMwh
ise1Iqmb3cuxuKtpTeSfiERsHL1hMQfklBAc07Zkoedr4Thu191PEqmKCFKQ8QkZ
mZDukpix7l68yY0ebHIFwxekRQ4Ecmw09+Aa2HxEHQzU5mqN9NfrAIv4ipvoROIu
ZQAC9HMHF48nRyc/OK9e9t4pP05g8yAaXnhpoiU0c8LI0PBbai3u5fhorBZaRcKq
oPRAWm0Aj0HaC11Gjv3gLdcrvzImDBzLn0fBy8D0OTNrCpNajnzxSshYwJDoeDHz
5scnjlnSwLUUxyoNpiH7nRik2w/MgEYG7+oS1bdawN4Z3PRVYvq0+KS9SD4ZQU5u
bU9OUhlmMwWLelyhwSVdEOOzfQWQwB4Bvg34sY0PMTdLQuUlZBb9yp03GcF+5P6k
CTGKkJDYTOx43rKoGhywS/sxtymB+6RnA9VWJ3n0n6mUjG0H0OFLr/RvabtMY7M7
OKrX8lIYl96kj5oivkj9Uu634odTKb6IXg3VggOy/myU0wD0BjTN9e0d8IaZF5Zl
5P3mXKNl65aFO/aNdcfQTgSCDIG5PZHVteRycmbsV/40HvH3gDvAKF8iQsh18VFZ
uou+4+kn3m3CIae+6gzvfSnKCi3sFq9lW81G9kxn2HhHzhI4B+b4NzVKHoYxKWUQ
aBSFh0puDJoMCF35IARFWOL9rPiqiBpd3fDwvfC5H7BR3CLJs4wpmfLFtiiRibtW
XI0IjtYVZw1GJGePfouUqzhgRbCbkpjfBKonCZefLEA3PmB5qIJIXPmPitZKn9F7
iVwywsclFSWqXYSpVSl2vV47XSrAaY/tuVILdE6h+/rtX448kdFMjG5mn4jvG9qj
q/kuuQVKCz/4PH3oh4Phw7jXVcr4UQLGo5LTMvKWWgUOceEktHjT3krXh+aMESPi
HhMwNNBgTv3OYkRUfBQTP77jmAyEiK3bg8jtZ9A2p+8nbB8xpBBI6eAt2tiCVAVI
66tT8y/C8aYH6kcFZkkEL8fc+6tbmu8Y1kz694nrepTgSpuuYn1r3oy+v3jSodBA
lRRE2uOrvqacfKq9Fit8Lm8sfFJ9X5HZKycXjlYZGHLuOzOH7koljrRTRLepiRQC
0g4s2Ae04KjA2oFLiylA7lmGrKAMOoYcwRkalr9zh7u1OrARbq8h0GUXzcJPAvbw
o8KxziSpII3LioswRqSFfFaZDZ+W8LmJisV+dtIyB66C3806tj8xscpee+htNrIE
ae/Cbim0H2Fhldpv5GS8/6hLFExysqOKRrbJXmdQ/kJL96RxlMrTIJobVP82VtGE
2Lg7hclNXxyGFB957fyia3uuIu8RJ4byR+gPgkQdstEKzU7Niq2Jm2xjSXG5PWNK
WMW9K9Nw6ja3LIwMRxeR1BbbMzopTLZcLfugdjPb5u0ZZL0AEa8gU8aWHqu+Q1My
yIUeCkshTNZg/umI16mCysPSR7tGooCD0n8lvMXVc9pYrEA8CRWC0Z5SNS/TSdxF
FT85ikBd7yS5FK9C4kOKWUV908EV0meBJHg/gl6FDa+aVU6PHxcTnBcqNL5ozG4w
76uej8GJWulhpkEtcrQs/1kW47Jqh7nLplyYFp85vWOA85nwHmDVwtgOtBt8UbCq
U7mFEzFGxRisfZ4se1GHlpd/c/YbCZAmIn5pAHhn9ogtsqOCGtw7NTe3sskVFzrO
Zba8ak+f4OdvlqBkEn9dMTXHueAHUpYVuIZQnva4bDQcXeHBjquzP4IY5/VxCi+1
b0tTf3RUVyGc/qIOza+PUjzAdkpXZvPvKCTSz9J/7xxr4C6UHD1hdxMBFFYOsmf6
wRm0llPaHzxPKAHAbxnr42b1N+i/pNpzAIbePTEaRjBoK6L5vkORzOvuT35GzjDD
OwiH+pY5sgJLobrN2Ot8U2h0zNcIvxtEnmYPUYEGn+L4NSmOzKD2rx85aENAUdLX
vPdp3G/w77C3PixMWZSrAlvZroIm0AZh4TO3/RS4HxNAmSnbf7XhwcTYVPjie6PG
DgbGJuW7Lb7TtZ1UdpX1qJ4MSH3Kt6jPMsuEW+liREsff59X3hnynKERoxCWop+N
ezTXW/Dy7Ie5Fdhjh1bXcbUoIzStjrSS8ej87YWOW2jqy44VrWl5OAem8DtEtOoO
iaJNyjAYBAwjRqM3y98KLN5tOLyoFAtTvFJGv0B6uDpFH4q1cvFQ4ACU6Xu8RYcI
9xoqpIRCkWbOEXdsGqQXqlvqDvZ2cvgckjpz4LydAhLDBNK31g+5zutRUqgt714X
D7iqd6s3cvKz4SjKTm2N6m5tf6oA4OxvJcO/4orPs9zGzG8TVlfM3nJ57Cwy98dq
f+1EWGQJFXVSnteazuiojLmWpSTG1qmAZkseRq3rQB9jL/R/sLzl0FOqGTXDHMge
P19SUwT+/Ivm8Z58f1bisvMyEJKhH0Lwjl/lzFaqJaYwTuBa+4AcBKtQoaHRBGeK
18EDZ01zq5zPoRwb9ogmQiI0YfXyQS9NWOrTjfql+ITVLtEyp02DGQZcOAVm4y68
gqCpFa9wYUFI72lXSTNduOcENGAjRjNIaSB+LKKvk1CGINSgbtqqD+6cYtziUZzB
nVujtKVSPiQGmhXJ4dsxkZ80VNre55HrWHx0o+pe9GKLq08DFVqP0EqkwqgOO+Do
CHmLHNuNapTsUsBZRgNGXb4sVVBEYu1J8KOTAJF6s3/TKo736VqXgqokcmgpJaAr
eZt+Fw9bLJN2ep6MTsrX2xS5xROFH+4r0ZKDt10KCOj/sVZcko4JZFn/icYx402R
2IlH1BpzAcid+L1cy4/j/XSk1TyfLrf9HD8HTcUaQxEl3Sl2tnnrCXebhnfv2AZ7
5JX/obSeJ+os8DIfTx74pq/J4qH1qjefMZF0jZedX2R0BrGk/6/GLWlHQdmsPXKh
WYc4Aw2iEL2waOPbNF6q4iIAl27pzJOkoHbHBB8rcUOPaL/sQG62VXTdVDu0dvyN
2eJSYWtnDXlopQdT+Dt68ZKjeyDBYUkR01IIt/dB5pq8JCaqZBq7lCime9vAM90H
t9fDkP1OA03E5VzOq8bNBSsTFt4CHRokDt+oaccxxZyPPp+LRjcHQPdiaZBbjvWt
h2A3N3y5tSOZCV8I3mbufu+pTLKZuSwKsp58gVQY9HxOMniGqKXjO/pf5H6VNKL5
JeInHJJT6vAyvc8yLNnipqk780/Rhamn4k0c58we/FvPnvDPYHV7OsI0KShPi/nB
vJ5HJRuPi3xRRE9MCByCSHX/5xWyZZhNY7XZEhj17wsO46BImGa1gh+FI9X+9Nv3
wwTdC4dxb9d5r0rmytHZWzymPgMBFFCQ40s7wc8y0XPkdl5RCDkhoB6XRHUOcGWc
aEVCRqNaRAUnSXaJ8IJz1jFL0yMulbkNjWB7DkVhqfg68f6x67w5e4uXSPaiKh1H
Sv8ffavIWwK6E2G16m/TAEAls1dWrAXm1AM7syIxhAbXTG7F/5OPL/b0FwxHOlcg
NmddKBEVGT2ewuyFe9UQCCDqN4uv2ytNUOzjN3tSbuc68JtYq+uurgrAF9ZLVWog
em6tP1GRWI+y7oqlwSwiArp9o0alx3oVK7tHpZhs74iWuTVB9FD23cdbUoPpai3c
0rvtcsULrRIj3XJmBUr09bpnyoMf+fQqQMOQAiav/R44Usj2eQ2zZ4GyVeWoGbqf
leB5zD1Tx11fNFx+1ke/uT9Vp09S/aBkrbLkkq08pSRRc7CUP0ilIQQnccKj0zVd
nPuQmM2Ih10PG5nYXG/LyB7i1Ibjl2HVjP1DSmXmFO/qIYb54fstH7urS6aM1ZhG
Pg9d4P9RfqtJAyoArxp8TNzpJc4QtZA/V4dx0ayH07vYmGnL/bK3DQxXBDT2RKKB
jU7nlTV2YuNjBhUuqQH8MHAuFsG+WBY/pQ5bL5u+zPAVukYhrVTHxxhsbRg144yT
2L41iBsqXXUFiNLH0xNskW9RTRciRj6Xut+d05pcJagcVZIQ8G4lpEIysu6v+N8c
nowsmpdzB1lbjtC8VgeCk+xGScPCXKYYV5MQW6eMxuO/kiBdFQOtP9IGTFnhUQVL
tAnXzEplj/vPt6pE2R4OBZWRfMZq7sfrz0hHRJYv2zK6/hYoZt9xlWQ5FnCb4rlq
K6BO39+iiwgtwT8LJsT8HtcrYKHeSlcxMhOVmDF4AH/tgdTYeFvSNvRxLZ4GHEXV
TyUS8qsqsscY1jDCptfU6uXuCFOvfPAvoqjw/oYouAFi2odcYr6mJeexRPZQaCsZ
sUO9ozqKxy9DI995LgkFwD6iXO2WIt51op1Jke+yO39yuu2TWFg+nSGXwRKBODNg
g0n+QxtbGq7uATTmhUsJ2pT27IM/KhDpE5RfZzLRT7S6g9Qp7P6HEfK1kzOnt1LX
z865inJnmJhZ190EFBX2BU+UAjRYspZ/o3LefCAXC9PT6gJxeI2rCmVPx7WGuYgf
jMblw2AjJA9w7dyPdiPM3gTGZwp9U/9ap0Tc0xQWqzCECU8DzLyvdawPAuMLGGiD
8NDsSvwulZmLdt0JBBX+zvrdL+H2IvFZ8sF/9eHl7NWCRjFomocMZtcoou9x0pLV
O2wsOUNEq1LeDrAmVdi+WET96WVWWQZGg8Xz8lb8Rv7mkiHFEtsN+z8J4ImM/YhJ
CEr38HqkW87E9pZB9xqbRDkqSZDNvEp9k6OSJqxbq8FkKDXgANM3tvgFBMGqvOmQ
TX5SMHVnM9meu8v7cj0ZDwRdfGzwOd6XuVH4xZoCzP8ZSzP1PyoQDCM3L4I4d0al
06gHcOvGYMmvDkb/rDPHwxABtNjK6T/XJz1+K97SFXMFjAtwlpEB4bSP94GNaA3+
WQ1SSJ6xDuYu9E58uvBPFCC+wqI5RbRuKFwXquvEdOXJROCpzHzmQFN3Q94VSvJb
XKYU2Td4ozYreb8gT/1hJf7F1TBZe40xZ7yPDKSl0AbuhGC7+WOsBBP01N4M/KLc
78hSUmuXejTes02vD5eYGZ322q7CVJfaz0U1nkVrGMtagemEU/sYuq4eCosBHkz6
g0Ip++HiPo7kfpcMDqsiPVMOOa4y6frsp2fn23BDLQMjhw2oyoTz4JwO1SVOohoS
iycg/8Ncao2Kyp2pmud5d5HEpYjS6+EkzNPbfU7LiJzIhuL8NvZcovt4RmyjA/4T
9CT3WG9w8cMOKRDurgaIXQsOOqt62rv9B9m2dj//uy12BX6LSzMgvp98kIvTEavW
bHNXbzJ5Qfm7lSJbIFeIViUgPnpJNpzo7jbI3KgpkBpMzyVqTq+z6Xb7kW3EHaHZ
pv3zfXUNNuCOv2w0OvaGIdDeL6siyHkvS6QUXitINyCn8HouWtvPbPWT40aYwdXR
QbyFgQiq4ZkvVbl90c26O4pojD67SAPah14+Jyjolk0mcjYAERvMoC1dglLT5LXU
WlXhVu3pWA/OqENjoMRa6GZaOqbus8iMToa7BpDNXPRGqHgMsH9Fo0KAoWWSDvJN
sfPkDPr3J38ETbs4W9ts88E7nBpRkD7A/w18+q6kK++C6PoGCWTfqiwrt5K1XScv
4PEAnSjxocPwh44N9iokqq9ig9DkftW+It1w5ts0ByqDHFKQ4WXJVDye+hWi8KKU
SdGKxINS8w7sr3fya8EuFEwpwnrLoinvYUfm5+eIXMU6+LJcdrRLGZHL1K4dsyP2
3L9bJf8jBpvFGG3qmOkN69camygx4tGDytmnfkndHsdulfj/QE31AV7PvhlRJe3/
Ya/b41Ja53O0XnsrMDqqs97NVum5Ct2NahpuGBOtrenfY6RtratoscKF9XSDXmxs
6UnbrdtWuu8hDvjGevSOtosnD7jP3GFfjV8/Z/IiWN3fD4ue3lCUI+pPkArMx9cF
zo6CWW2cjzTN1FpRax3SzWnJyALPVZ0+oB2uXRXTJI80Yv1KJrtTpWzbWuiFHVLC
M1TTuBLE8lrlmSiCfsGih67WvKlGyxLdSpuovZhhDqTU1SknHtqWfkJOVe8hrUFn
ckvkEU1fxsDRZdRn15penrPN91iZfrGwkEHgGNJ9MZlfosxyhdnhh3xPFJikL4iw
aeqVcw7kPQkTE5zGRUOD+zScWcwNNRd20X1jWzceQ0NMwBdvYP315ZSn4hq01BvW
Qvv5sGabJHjYWmTAdgAxUCZVhG2/ofmJRMiXuS5EaSp5Bc6+U/G/3dAA6XifYU3/
uMPVUDR6+PItj85ZXAl9Va6+L6+XFLW1rCGNCcXo6uY1kKbOxhGL1Ms2PgUNlT9t
5OK5oUFbXFGjjgXrGFJF3oYi7XwYDdISYmxIycwyEyd9gnvGsgLqSHt99+Bz03XY
T+/AweHZfzgbqdFNx88tKxqolavigOMJk+SHFTHaoevJkNFze5uwKkfEcYMT7XUA
en+wsVLV3HY9U37h2N5iSM62SZqAtcunewm/zC7lo0VJdURnSBPXaZ9afsSBeLJH
+4vxl4Iyxriab5swKqki8mCYtvZAHSY72Tj3YoN6rLujn1JG/LijlwJS363iNkjs
CA+JmW8Y+cNPT+32/Uwap6bXJEo2loNli7xiTfdK7R0bXicNSbpg0XSu6DWmvkCH
ZT2hxfDaNlzyTWfsm+R3bRKdSIEgUhCdf+KdFTXRlhRnV5kU893QTXotc5vd3W8h
BFQxVri4upUlWwCElZuUUpUucb208jZyPLnYZaOOudzhS3MXZwbXDY9E5SG+LzHk
/gRRSc+Y/gaykK5aE7MYYFi/hNUDwXcshl465TZpquzfM/t6fhNgQr35WzPbsXXZ
lhRDGBjJX74emwfC+rKf3KrgE+IOB2JSsbFkpCNtxyPGQZVlb55UXWbSDdTiZstM
3dsp+wy3aLe4qAW5TpDugzJW7yE6NA/zAFH04IBPZyuvPyDm8AwuU2e+d95/Nn2F
kw2fqtHYnOzmK77aYrW1Kz5HkaKX4LyYVvfdOmk1KCp+SoQsfYZ08Mt3DS4F5Yfe
XXSO5kJidlxzMHwbguF7e2rba1A5/L9MaG35LPFvIi4Fspn6s+CLzGL/3LUf91oN
oR004SwCtig32bjWuD5rJoceoIpELVg3BwsucxiVR48WrGty3S1dGiZwh2LHenns
eNZo8/0trkDNAMeGKgtcZcHnNlaDTnUp35wVe31Su7ZnFhrjaZsOyb+6rYKx7ueY
YX8Ee6oNeq7PJgRCyPhfNLU9xTisfzTQgsxZHEKr1SaR4YLBmArzXL72Ls7RDH6T
Fz8UFov2pitvx9MiGK8sHu8hltLZ3zlO3WvoBerrC6whvGAVgJHWBUJRXSSkpp1p
po3cI41OQWLAUE2lariyPDybUiWWVpbv6t8IcfCiFbqCBt2fnkYObVqQn5aZPw4k
0jtSGm3fAPxG4d8J1kW3T1X0Puc1I/I+yjWwNtdvATFPAX0s9DUpDcFH6fwNoTcx
SWn7AcamNDBUm5uCDriZ6G/ob8XUinYXcrFLFYH4qTAo50gFodeZ5EDiaUFHTIdO
dDa4SvyvfL6zNQRb9OgZGW4pPgollWcTNUFOl2EL6Z83i3OSWV9JmuEdhNz5LfI6
YO8FbRrFBlG9+npdTmyGcFi/9010PoZf910OUfvgmebAinMEY7Rmx6+MqSDNcX57
KDixkgFCsgOeuc8yunMhv/Vmllaft+gGNf+7NrutqYUw8AenuHi5ZdzikS0LDGqd
4B2IGw9mu3kaUYOyJIaEzCoNvgK/SpA0GkvaCQkRQkdC0nztlcbMADI+54r/yQqm
RbNeuPbwCc59arffDBOisAD4IhZPcmYPREF9QMuXIq23jd3oZc8hqqMQ5RR992pD
pSqvBSDS1NhbjzRVfdRD3H9B74wADP1InzmXftJa1CuhEMTA2ZzEuskHtTq5GooX
EaaFW5nREmUGE9vHO6fOD0if45/VXbQPVn3EWy6bnBzxGFwmDqoB38A8TaN0LcU6
479IQ7oNgaU2yE3tcEm8paNKtJcvj3M+Tei1wWi2JZM2IMzv3iJGLRXPjrT1Vfns
dope3MHQncCGPK3/W2LrdI9SzCu7fv3v624RBgysWwThg/mkKALJNZgMQVZGCyQ1
NJXV+8twTw3z6EWLB7WaByjJ6F3ZqBIvAWE2F9KJSZ9EArYCDHlI3z7W1eYulyqE
D+Y9I1u0lrOp7Lp5lOxuQmh+IImjXsRFIpY3KGSAfSzWjsBk4/t9omIntiTqHMan
0mpjKxJz/azl/q45ul2W9dJWI717Fc2ezFy8bR5N5Lsmm28ez0yyIDB+vei+APbW
CTzAsEQLZKITn5rdWxbrTFEY2yle39z64s/MTfSbK7uQ4TClQdmJHGPEaOsMAGbU
HRF9UIqoWxfxui7QxPPHeZZBBmyIZ7mJWzoWwFA+hat+Hx/5X8+KkzWbKneBeP8n
TRdPA0cwgnFITxHXG2AGWSyQkoQqAtQAaeIWt72v5BOU+hmBvOa5lVXe24GrmSy1
JgdLJGnpmeVaSKieJqUgkteuHfXmNfn+R49vt/22mXS5wwHjesqlTMCFF4obY+bT
gh63WkyccfxE3/TZZh4vNM2mwJWFR38EHu977KPA1eW0qLZBEYqG5dR6KEtELU/V
tE+sRTQEmYIHdVv8CjC1daNWnzeQzzoH76xYIGlSq49FYLjk6y6u19608U+EP2sp
REqigKIhCacjUg4qLoQrs2qASeJJlg+L5iHEh5vzj96QTn+ECycYx7GeNozI/g/D
IzELq8FBYiCNoST8beTrXopKo+Lon7YrjUKw3it06f9Ja5yVWd480f24lNmLec6d
Ik4XEMpZwJJRVEdxfQvscfWF1QIXpXSPy04gzk9ZekpBVgiId8csCmJ7ZPGLxeXr
D99R2IwrYMwUVulyqfVmnmkINi9MtYLP7M2+RpG7j9A1ZIKULWo7XmR9YXVgaBWh
Lf9oY4hb13fmbEX2d9YyZh5NUW8M78385VwYi1OmIvi0JSkAkUfM8JRyxdrUml7+
dHqu1IHa7F9v7vTj4R4XduR68qiYeLbtR67hebb+NW7yDnIk7MvxfD8/VjJRpACr
fp0C9R6QEFTzWKp50qe2beZ+DXNGuFNC8yX0NTcPjKQPQ7CACvMKG/PIKTA5rAzD
kAE58FEas9pap5r75IBZZbH/sDnSwtXDGwPZE8J+C8L1su+nOsb7XzP4Ign8Jdw7
lRzWm7bqs+y8j661dYbQCm1aHC/L4UNTSMuq8axO4B0c0HIEMTHseI2XvtnQdQL/
44yl+bt5czd2so8wQ2Qnk5aVZpG3ylImxjRiWmn6UoF2ctwOKd7Xtx0ZDx+HKjVW
kO6JYis2kkLNwwSfChE0zQgf9mqRVaEVs3Str4KZIqlHfNwuKbfyqIET48i4fvIb
i1sBn1mlbORQQXG2lElR0v6uShDmEJwuFlgPOOZn+HSdX8CbGvr4EepeLG8cTY80
H6feAwB7tuRUUX3oNIs/Z+LgknbYjfeS6nTPwXnhm3MeWdIWOwrfrSmkDOn8TJk7
h0wBGd1m0uHkc6POf3rrvMU9pF1sdVI8uH3TiXKvfB//oWtV0IX1umAEoja8AWHm
fHAw1+neMqdAz9ik5Wq+lVszEm+fzcbsuk1d0I3f6AYKxnD5o4LAirQnaPzp+kS9
Bsm9qLscJ36/aAdzIFf+1YPGsbk+DRqkCsfdZ1PUDUMa2fMGdyZ1DWaoah1vprYt
bxUKOPKDUqBug5qYYfg0xmd98J6TMHs3Kn0bjOw5EVXXFhXRm5OnN018W+1yjjRj
BCHo6pe2p82o4Rf3DsPQNBVzlYIoqgGjM25t68Z8hTf5uFpEbK1iYtPrKZ9/zVmi
wnZt24Q8AFc/0XorMj5PHn7o2JXoQ+4AibXn87rVbkUJ70AjwUR8OCHj0TwLdG/V
PXy3cdemLujBg6IuqisDCbgI/kMNUXMWrZ8NVdv7YXlLIlOLjerSV8/3tEHNcIA+
5OICopCaAHhm0tXVl5lf+NTY99A8uMBGWyd5aXP9VViZQrtmwTf3gTxsS6wSKcYD
//pragma protect end_data_block
//pragma protect digest_block
KnUt5QRorHrP+OPQse0f6H95rTQ=
//pragma protect end_digest_block
//pragma protect end_protected
