`include "Usertype_FD.sv"

program automatic PATTERN_bridge(input clk, INF.PATTERN_bridge inf);
import usertype::*;

parameter DRAM_p_r = "../00_TESTBED/DRAM/dram.dat";
logic [7:0] golden_DRAM [65536+256*8-1 : 65536];
logic [16:0] addr;
logic [63:0] golden_ans;
integer patnumber = 200*10000;
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
txTCSQZJtNwTCq0J3jn/9cI0/n+Z28SJUdUfeojWpFvj54zZvrXTFtAluUbao/M4
QPLqbK2u7wLjK/aLKMC/IGz5IK7Bvc2FZf6etn41dldeYx9eEnO/lpa0I9CY0mtR
ztrQZIbGsBM9/CFqMo2jzvUiJDiV7989M7WV8qIir2E4XgFLIpt0qA==
//pragma protect end_key_block
//pragma protect digest_block
AuwJsgAp1viIl3+/XviqTnt6yTc=
//pragma protect end_digest_block
//pragma protect data_block
PGIg136bY7+hGMERqb1kMdLNjk+7X4Ybv1wTeYEuG/7CmS0ozJ1dwL5Ff/a847R7
KtMXtQBm5xBfAnhvOPsDx+8c9LSwAEg3n5OjgqdM/tORXff7ILyykR6hL83oc8D4
M8b0AtH0pgd1iLgxn77gqStoXvspqPLLtwH6SZz8r5FnUvv+zSxgQ9P5tFs5GwUR
9cdbeSN43pDA4jr1uURn1dO1FfPJkcRwYGe+Oxp4Nc/PUwwK+pTzxHMoe0nO8nCa
6npekJn5CUoG4tvs/kb1wabvyRnpmRK09hasoUrhbD/CRafMCzOlxHj9ZPCNlunS
rFEOIpQ/skrxt0u3v+5pYsAGCNsrh30zbsKNfgt+cdjX25F/qMYSGzcL1GvYVXfz
FIJ50gTGRLZcMmTXOoMr0BDON5fq9KIFXvJ3uQjFYzNuXVvMok7ThGOgvVsFVtcx
KUGggeyzIqm4eYjz7dsJACZpeMCW/1mk+s5yToGz/mN61+QV4WSmfgrtOlFKNK7z
fN69lI3Qe+GtnBnQqRd+E6bv6VdxfYuJ5bUbVzWX6sra4qPwPb2wbQp2k/zSgo5F
oD9k0oOtwfD0y1hxJm79n73CrGdS+sKqLO4AZULyDApqKXFlIqOR3UQPi38elLtG
75qeBL7QFqdbAtFMJSfiAqci8AdK7nglWXr6gABcwG3DM86/n3Zvm5od6REbwXSm
pwDFobyIV0VMabEDaF87MrMjjYSsOSQdzhT1kDaoplBIBlBmcfdopaLdp7W+2ouG
63db5T4oGuIC7wUyfCPkTiAiGao/poWznFNSmXAwwilWp1t0YQLnUulVx5FUCZ/G
KLWr6ADdhUdAhcqabjCt0FAJmmd1cVQ5y6tA5g7h/wuZ5Fn6rrVXUHVMUOEEAV6c
m1oL5jeZh9Z1hN9gBhJKZS1t3YO3NzUZOMHOAwMGU4cjIKB0Vdm/zz0R3N5hJ76K
ptCIybI9t9YorL+zF5maPhfSAD7GFfgc8Z9v9twGS85YA/Pt+iPdg8wqiGpyEwjq
/b+vKpe4xOY8PUXQpPEVDCXddI7qa0/4viBvniTSICyMEFJ5WVaZQRL0yhnIKkn9
E6YOWPjDq/S5vxqjY8vOU/N0dxzhIUEnN6K3N6cnpwblw6H5fIFmfasRIadMf5AW
/1i25IBAeKIjHyOrmDx7w8eU5ToJK+PrbyJvV17yNyyz6bgHTON67KXJfb4ygHJV
DN60zovnMvpn3tnQh8u5WHwYeFLNU17BexHc0aF7b275uHtJkCSuk7w/Xj+vd5ze
KPX3o3JeToYLn29w0lck1UwXxeehsMkXFBU394Lk/JQ7qMqVejUItQzElW4zJSGP
S2NjYSbo9MFtaCnJkhcGeHSYpdWuW1KutmhyCKx7JLkI/5nOLDYAQ3x1sStXtMli
R8mtnx3O1FcKctpdEzl2MA7WVO450+Vi1FVfRAiP8KABw3GiqUL1zzp9kiErhuUY
KGQi8UX689Dti80VDGu21iW/lSsBHiA2Iu2DGViIeE20Syga5+Z++3qvekkac/n5
vxoj5GpuGjJ9r4cNW/7xh4ZJhvBcnDfUTAXDq5LQmHvKw+5ztGP0uP5T7fd0jO68
jqaJmZ0AC6riIblUtJVB5v9YVj3tk4Qt0bN2zWUV6JRWQ/kuSI+fSQTXeI+7TDOM
jfOt3J+7ejMojv2nUEAKfpzsa6738GjdTvkv3s1rNe03od0oRYQ6wmb0WJbOCJZu
/QHadefL7fJcNYgXx9NTUghvFMGgFs0XdSIxjRyVjZd9fPkdPqnMRY5g5b1oubPR
oDb3LsWa8le6avyCaTvSjgG/0OAousJD925xmM7QaTrvWkqbtGycZg1Bg2fQobc7
M6xZDdME5YY8tBD5LcvuNGCpcsmTCcKQOMtOFi+auQdJhFYmaizXM3CaVzTcGBEn
1+szhTmEgc6RZazX7yiVFS5EmIlDuT0Epvc8B76Car26IBK4XfrzJHXuCLOvBaWo
fFUCAKbgQq0KjOtwwjRDUwmw4/qZ2ng/IgaQm8zwwf5DFqvbXq+Z+HDOQvaqPbGg
nsJXG8IMwlV9jCrNgT3lblgreaCh+K6rWE/TZweh1L77lnWCU0GXxCVxuXFH19pH
kLk5nO1azuvglHrmnNGa0wJlAdVCiLSsGssB9tLmh8IfwffNUP0rd0qG97mi6hLs
uO47U6/1m2RGVzp0Zz0bSEosiRP5HDCysMRT9RwgHwBoA+g/XNahHglniIN9oGFI
40XhhjbEe3DBKh4L8GoFiOBzL+GLFpT2fRVlT3/pQXavU0k7Pr4OwmJ0PqHw6T9i
cWFkrDJ0ASCGi90QEQXYPr/IRZ4EV2+hI1C+883kUgOKeWQF/5MmdIAXB3kJTZhk
pDpsEMLSPaaEXYayYNFWhrTK89/+qAidieNfP6A0Az73Ng7AIiv+6eRvAdzhxGbY
zHH1MAuiA2EeaoNGJ9ZC4z5ITtJgAYaDyyBaiMqns3uY/bwRN5Oiu73he3Gc+xUd
on4fT0SDEb4q1eW/8vf4sGt6njsyO1025ILGOLoI+WUgwgICHkjIkafiaDZgflGM
/AMe9ZxtkIywX8uTpIc+E12wyD0nq8pbgFWeqOC6uzFCsopz9u9YCXeHs+GNEu7B
TXGnCD5NApN3rC7iNIl7I6Wfwi7ehC1r87KfLbdy/o39H5TqHW6HpbG5EeB45uqo
lCkPGV4gpglP9H7lgT5qdXjEIjvQxPhljBTuwX2FqMABsM4ji63j5BO9J29d5oUk
RfWOs6vtCvra3fcZCSPUjWGOe+N+LiZoTZPA6WQv6gSXSCAnzK838sFXnZnt3pG1
iHxN/kpWixv42jVi8MxFGzAfq/B1boL/3XBrrpTLaXRt6Lu5sn+woKQlx2BGGrUz
db9RE8+QIOminQkPtWsLtc2l8EGNZGtTPLHLD2wIqIO+CsgFj+Osfzy66QSflrVu
bfkHhSRs6bKBEXxGmn9jam8CrWpQznLFJtbipnetTxi6C49CpjqV7exC7afcJaE9
u1MfBKS5aGjtSZ2Ka9Cc4+Yx3g6tP2Km2RQDYYKmdDBdGTcttxUrO9+iywl5VQWV
RrffZucOF2C0p5KT0u+OWtWwVgohxBjsKgE7Hq2KPjV9p3249nZOgzCVqIaz15vZ
6JWdeWoW7FwAlyVSdVaLQD2atEk4BzBj/vSHLQwGNERYnRgOYwzOePzgNj3H38I2
/myV40ALc47fO02Wiww9bg9iGBkS38U8GQZ/x24V2Jx6mK0PxZTl0nBp8odps4KG
8aWY0663VYUUnYGx3th+yC0bbeP4EZTLKsl/9ZgxT4gtdY/qwwJKTMONtmXrq8zG
Y+p75QscyX2zSiCKJkNXwRWjATk4xnXDvtN3Buq89dBKz73JScP9JUFBKr9Gwk3L
ZDqOg8657lB7XpHxA/ka7EyOvdwwhd3O/XD9jc7y5KLxwfFEqbU849XiG1zLdfbZ
U731mOXFInKm68dTyEVBvJfdvbzOIj601st9ec0qm/PcI5hDa6C835AUIhFraafQ
osFsmHaYsUx3xg9QA7sSBf4DpAVPfSyqyRRprSSM1R2B1fBqCqX/xEi4uKOJ27kq
/OunZhAeHtHOCvUICZzyoMTJbdWrlDoKOc+2a4P5hKHJcWKuDt4nnYmauhEA0h4c
/uYb7YXLQsvoKUtJ8aLgyyS9UFSDqdZ73BIhAsz6NpfYKG670eQHKVuF0ZvpnX8N
mZYTxkNBvm0fr4RdZMd9CqvWixafqCt8viEJ680T1LRnZPt7/zS0mKXsDCmMvYN4
G4H6G8XfxFlgVMoXIVJoqo5KK8JW5BxzbsJzFQDmMojBKxCovbfogUAFRjneGZc6
/ZBp1leY6f3FxjqBOxYhb0zd5OnIwUE0WWEuas99ImnXfPmP34qJkHDJ3H4Fg9Nm
TAIeX8ALWKwEPhSQ2uQ7beC16a+l1E00NOmuxRbUas5vNGvB1KV9yhjMhYdVxC5x
GI3kL+B4I/Ngzd5fZPuRHkwQ08QOEHUbhH3eYUm8TA8cvlLPmY/vy2B3QrvbmFC8
9/2BlUhLuD+hQ50Tdkv6b+xwTttSWipGD9JC2SatYeRdpvY2XRiUYaDsIvC/rOR5
eBkc1G+zRvZU42lqN0nX5AR/J35orYBiYe2MjegsTU0HtZp0EVEZK2Dj/ypGnxu6
7eVDHiVqMa1b5TiVQl5nvnAyJZYOpSSyRkOjGOhT7zXuyLcW5TeFlQqUDIXZTJL3
E85Xu3nfz76FQu6kjMGL156tO3owv1F6qTFaD4mB83SlNWJ2e/1ol4t2T9dzMGcB
XoAhks/XhBmseAwQ+9JtUPEubk6fJdpIAMjgelqx92SOt0jEmxMcCUXwT/UBpGF/
UYpEjrkHLtHWcSybWjNpgCQ+MyJho2P+K27yNYHrrLPsHLrDqyq0w0nH6McEXXxg
uxuhmlyWF8Wx9eFsYsQO1UtMKOIamszgMuYbkgiI78UfLePAhsOuxgcNORRcDIbx
hWsyq2kmpLlrUDJDBDlmzo42UKRXzsL+OJAOknpYBLs0CZ3FjTdeIOSETzhtv9Or
2uFHvL/WjdXxLTkBmA27CtYafhJAx6nF+hnv+1xkPKynKmDr5eBCMVASM9wWG2rc
QaGU76ZUSYxy53/0rCPzl9iqt2KgN306vhxHeD1+EQ2nXeF1QCF8RtcQy6hQuf4U
iurquLMKXlRA/hirZ3Vj2dSNl8YTxbcp7clHsfB1CBKKZDWRzrrBn8CnT9+44fjl
6eCW5J1+Q9vubNpjyGo492o/j/5IJXU5AAAOlRkJaikJMRyofsz0+gWHWqJApyTP
mZu2m8NV+3xQgNRavGfAzPhKwwpMfHUcYFwcwmDoTMERTZ/0RCAyuH6HMf5DWIPL
/ht2NLjsPpTqogLVSlPkH2Kb/TbuKdyaGVAeElUF5rB8TXB8ek9VW5OyiS2ggWep
BBRKoJGvbqQMqdrtBe0RGPa/scRF1kqh9xc5nT6c13VhUbGI9ojkQk0E95bdArHv
Ufci99LsSTMqWcHABIFRHsD33zDCku5UEKxinNFy05ZS4gZkMudjU9N8Gry/SUap
T1weGCObTU7mvAQJyesgyx6f8dUO2wFU3pMY6v7t6lPaxd1/ywQ0fLUtGppBPgn9
FGSKU+NYQ2IwL9I1ma29j/4smUqQRNTz2D16uRHJAwdJa6MdhMjCqJdVyD80B5pN
xx96f3gd4XftrcWQ4iWmioPytCnJToRfUnMJLdwJeJEhZ30rKWxDXFjHepelfzys
XlCqh8mGfVLlvRoitC/eYlIztPwCfDjC1vCbCoy42/3vrCy2xt9Zx0bU6ng00Wje
o9sB5rkx91rcLLJDMzw5yKTxjfN+8ZgWB3GhderZ7h1sBe4KQW2UGrV9d/yp6LcU
IDFoOfbFFX9i3rSm4oRk0x4nWC+uV+NyA+qJ9na75KOUtJEHRfaldaYeAD9NlfTm
KSPV6y3EH9olknx/PNGmX60o0ovfqI2hVZNS7Eq9UFw9YOAqXlAw4vLAk5TAfFuE
0MbcCc8wJqZH0P6HSFdp+LfvlEauZl+WrbezqoBR/PfwOOGQl1srQXeBEnf0mvHT
WlstmQUQtp0kXn6B/SB6PaeBNZwMIJbWlh0XDPnJvqaxp/kzOXvBaBGMEfPd/xow
D1SZLwCbUEuemSyD51HN8jbLTp2iKJv1FMarSCXGIiufaE2ktcoiysU9QIWEPe9r
oP6z4gVVaTuZG+KV8Ml0bC4AqfUVeve9AvN21Jijbk0QebK4dYGEqN7VAL+dCwIO
T3b+GHS5fihD2qUtWW9FKVU9hfH8nyGlRmXi32hiKEvmKpqIKEfZJD2EOduqT4yv
1j/CWJiS0nUYVlH8YhoDkgDKfN14WrkVYREaNgH0NryXlBczM4MsFE9V17EVgkEO
VosW5y1LnSBS8DvnieY0grsi0jSVWuwqN7voix4UfvPIZvhThf9f0dBeY7gUqnKX
YoczeQsSJ7twKKSOy56KkoOortwSBiKcZlh5ltlZS1NLq1AaaIEGNaSFytub1l7z
Xn5GbolHfHdXhsX/1Bj03UOutsFAfTczobcAFKATuS1Zi/DtGNiL8MadHEqr1JyS
B3KcijIJfr1Lkg58m5D5H4FvGsDoq5jg4jltvBWx/mJupfrVF4YgiW80D/7StGu4
7NEhMit92F5zcYP3DsFCc1S1XKCvXPzcJML8dnenTR8KRTanJlUQDQ3idGSJUIPH
FN12p1fzrn6lOwVsnn0tNGnB6FricukYjOwAZitARY+f3zi5YtbxLQWJ2Bhn3X6R
s/LFtqpUkLD1tcxmct3TBnRBKdO9K+sxQHSVevRFnVBfU1roOG/fAhG/DI4odRxT
UxsH69jwo9xuKndeAzvikHv4xjD46MXP1l1NTzwhIGocSsmmT31a9iqK6Wn+tL52
cyJVQdveNHywUa36SwCqmEt4fZSfNxoWgy7H05MaS05UdR0x8y0VjiCajkxqaUhD
poWh4r9RsEdX7fv/ki0/Hyzst3YpQ7uGataipP63YQbYAEa6h5sj++JizGSmdHt1
sxfdJRd9D5nagfL1LL0OaZicIiyyxDry7232549qyCE0OkdsIYa9EDaJmV0Q1igD
lN2GpR59fnukW7tphkGG6C50uefSeIiV+MZtL6M3qPdRr4EDeR3cNMTD1zqM8Gsd
5+nkRTmQA1OPJO0QpyA+tjKQXpjvnm7ITLBfeyXQXUmbqRAu5jyFgiVDGzU+z9UF
/6GKjA7hNZ7fWJUUGVVn1pacvnj6rNIQ9dYgvoc+XDH+/ozxaUJmBLZYz3i5TlG3
+sH9N5fw+m5x8hZopSCoqzPhbDJ4DkDGc2ToXDH/FE4GKnUOgoLOitu3bWtgYoDe
6bCVnQx/fomRql66RphYFTEKx874wMU5ILE0Vf/ADh2lEg8hl/UJ2yEeGJwlxGvC
5awswxJp+3KkGQxKLe7FmTr0VUrD9zLHetzJXViNwdJbjTlWuLKPVezrw+vuHAXh
gtVef5GMTGirUYsAzE5zTAn9Get1PCG2eUbj4DC8XzalrwMrKBN9wk8wu6x23xhL
uBL3Z2TyWzfv5uiPUNxMpvXRyCb1r/NJPcRCMxz2IWchdy2JNfrypa/xQqPlqp1X
2SHk6Nf1G19vVBgFotlffBFEy1FlKTSr7TBLbUxA+8p66aAHdPrMsjm/x2QKJoJi
ZbLm1rX9EXX8s8FILhr9lXUtcOdW/a2FG8NRayJRLOM5gTULeoZEuPZAJHJ4mNT5
3gB5XPwUCwAuBIGNYy2c48vrsyKl/Nq0LS2PVW6qtdl3nj2TsscttDqza9MwcDag
pm7doi/FwylrSfr7wzrLxe8lHLO42i/KHenZTPh38MX+GfhsRXbxU+hRsuYucggg
aKbkcCzeBneVkV91xqa/hEgg+CAfxoUTJS79Mfykoay5b/rx1dMJyM8e+yI2fjD3
n/WYtlYtkiWHt219gtUfzTedyJxID/aV/A0nMOgkBTdl19uOj0X8hIEpZ/eyslS2
/D3C0uu+YBqgfBTO+pQfoXTiAx8EuqpINjzKJOvz2hm3qdzZI1pKpr50sRX2YdkS
7SCKshWEtZhrDb8E/+tV0c8MTlXJ1Xh8w3x0ti34B4/ej031fPpC0C+dUzLPUy3/
wvn5fmqq50CzPHOhmb4EKPO1taJEhc4RWN0SdfBY7ZknoUq3GysIVypMXb6vfvd9
niTcZ+Qk9ZVfx+A458avLWS6AyO1113E7TEG9ScQeF2TmuWfVILqL20Co5HDBEMc
82WKZaZeambpBjd7yx8w8tsGAAfAojrJkf9JZqkRHOeWVDxBIarFXLkA76Qvm40c
hrIqzK6djm/tZiXFRyqqdcYOmn+MfRx8wqEKEAcwZgQf1XR4yHOylvj0W8W9SCWi
gyAmK2/TwAcscWEOzoqbMMz1UH1ZVINl3GlFdPThBduWLsJ+gpVzBt1nOUi7MhFM
yuC57UXfbvBznZHtC+5hrDvhL1Mp5yfRfHu0mNvZEmn7n5jVSBLng7lovc9I4Hnf
Xv5FtyU1RSLF3/Itmj0gFCdH0+y8Gz2ub9CVxWkNK1Wa0hA5dm7GNAvx9e0pHQDk
FbouEsrqZRJW+1kllW0ITFZtFs2z3rdQTKsB5NIptEi056RfNlXnO/Oj2vNtP669
12SYG/7XGW5ZOPW+WtixhyZOoBxviIHJvKLONF+oqIn+PASrXrnmBb27F6YAiPH6
THoBw7Ic3hbaIr8uX8gO9jykrsV3+OJl/VNudAkaJOiD3Ju0fiizzmhgAV5E53/h
1MA9aw0rw8YV7lbQmOxKZ6G85k8/RYD4gsxBfyv/6OCffD7my/IA7Qj1ln41DnQr
tmnSdrRgDBETu3pgviyEXD0JHbnNVgpyvZsPiyX//fHg3FQN4A1TT1RBb0jZ5xFC
R94q4OUg3gGFjDe7lu2BcDhK8uW+93zjvRv1cXeoZL11z8DNwk38QCqbu88CqrMZ
bIPH+7DpVURX4LOhK1wfpCRYgKqTSVbiaeD6rZ+lRYiXAZmzBquxJPD9Bjufekiw
qntAvHX95QlbFB+YGyXHZoaQSszTkmicKS73aT+K6GpQwDEmtGXKa8qOp2ZuxnXJ
xbXmD46hJtTwvOr5/Fx2k1MqfyJKRHm5GgzYaVIVpWVaj7lCAWGy5KI+8555YKky
oyJqfVNACDC+nFdypuqYwkiM/0286GBaEVgcROLu2EQnAyz4PBKIQE8b4CmqxyBG
XOkoesLUSmCvMpc9tJpRPRGom8pQd4sd5zESa52RaJVy0kqE6hTcn2+GBTbj4Xtx
SWKeNdWHMlTPmjVIbBYSMrvWrVQS9FaV1t104z/yo05FqBW8+esd/bBq1p1SW++E
zqLYpqABGVsDu5/PS5yggANPFNpcJ4sihunv5m5QOjZnhhb/JOFT6GwnulV2zXhp
bfqL4tLZ/PWTEm/yie1qJfIivS02im7alByMad+3ryKHdFDVOJI+DDN9VEw7wgi/
UMI0WLGY5ATgegikim6rICVaWlSaMfQ07PHBc24zzBea3kyZJyr9iB59Enwn/xaB
ihqz1+CGWNoYonprjDnEajbaiJaP85KoHsS8yKEhvMvkkrv2NqKIvcugHCPA8OVq
8ecOp6WWnBWsyKmf1kCDOG4gshhWDEKf/F0hBiFtw8WXeFTExDj1Pc88s+ws23+2
zc+CAuMfxTkyQwbG7SK274YkqeEZmdzAXD2G4JJ5xcFvdd4O9o3SSNhI+kQlyRQx
hXsJJuwH+B7MzH8E3V3AW9XN1RC4GKCzNxDtRLuhhOBXhPS0N//8Pj2oSIEepiTt
9oCejny4gAwyJxXvPQF8z3Zifv4I/WBCctsYyTbJMghtBZ1qaEtwJStVBEsbz6kW
DMGsRL4hnz0+B6qs76imm7WY3Jrt/U3AVIve6ry575+zVQwygbVM7kpsgR03TiJs
cHcHRsQ10+fQgIAFwTxODZeuuh3eejqkPbDvvVfNF+7BUqaBlWgYZNKn7FeNk0Ly
aIniTtFs7hgnt2G+JFkkIfO27SKPJCVhztp/+dieQP2oKMx9+goeMTnijA79ZLiL
S6ZasI7y3X2Ts+0XkPyMH0DMZVD8cKAXiqx/eyBLFYialYwwYo8QtkDbXklf44+7
nCXIw8fpTrN2he24Y93DODVknE9APTV/NkO2kouxEl2ZcMJCCzvLWXuG3wml128W
t+2HDpHkeRg7dQ0E+L3iQ9PYrj2AAXOuGLV0w7cPbGMgkjEtsDx2Y/VMx7tN3rhQ
7pOO3QDy8acwxP3ifkfsoPR0ywsY4rN4p6koXqqjWhielcS9izzIKeXc2hYXW1Z3
B2k+eV/fcwtIStRbpq87Ac1WtncBFgN2pFu+UKYzOWqkaWIxlHCBL511gcMrHAUS
m8oU3S9th/MKfHeBmIHbMHbjUeQucEJT3n0xye2Ctn/wJc7RF5GE8nbM7Izjxci3
F+WTMgC5CL3NLFHPR/EMsvaM/lAKsfNU/pVNZ7zDQSIPd+rAj6YcVkFcRiREpLgY
9xEqIpWHMSL8aiUaygpK6pB1arYyU83dAoOWfGJyUMV58sjrPgdaigvPdfCno1+O
qc6xICUiHebONdyon4t3e6t8rGMXnUVOSIUBMUTMga9sB4M5SPVmpRvXCeC8ssxe
0zGN9l6yi0M34g8kz+xsn8XvhgcKTh0fpu9Ee/hBUMrDw2av15S/zoDGF29E4xDs
rq3jdUY6r65NLY5hb4gz9wQYfWNsDWo9tqb2GITohr0vFdBD9WRA0epHtUrZ5FfG
BbD3jB7wzkbKE5TU1PNglea/W1AGW1NxPtUgfkdtlQq/Xb/Tr0ogDldmtbK+Ur8d
q+1GgAznJHlYQnHBGb0bxfPsffQZ4SQQngbhfQzfYfHloQJUV/WS3VoSTI6+E9up
++GzLU38sMJgc4RJtaDNgjx0QMnnyYGFJRrgtKKmna/IzPHPuTSYvc8P8QGY5/5F
r0R9oTwdobriImYOo3RDtFoJlTK2QOyu7QLLiAzJpm2uCGkfNZVG9hGWtIwrrMNa
Dg2/v740RhOalRToKe2m4tkcusl6SGkWXTA3eGwh500RhA419OOH49v/GEZYo/Nc
j+e80DbNhT2Y1omSMCVOSbbc8WB3ut73DP7ZgDGT+MpxdDjctQx84QVQHRPDm3hg
II3aFzuoD3GlpclPYwUtvFYaq4jrCCs4Y8OZlcNV7WomY4PjKYOnhez10kk53RSy
kxRpz79fstjx7LanjtxRE/sONxR7v1U84DqC0/EL0RWXS9Zd1Lzldvq/BvzFm+s6
p0uWCYHfi5LCcsHgiAObdhUKrC/suZcYxthNw/6AeddwlakgkAW9asxLKpOMHDhy
diMy12Od4tU6sJfTgZ+EBns9YpSyD4KgLk/L72hsPiY/Hj6WJVbVnQmnKQqR44eL
bttYZuGqr49UueKGc6mI24vZNFxV8HTt5MFkEh/ROawRqFFBob+aodQwvjqMcejl
UjQA0DEjFvQJ99GqLiI4sgb+DJDE0QIdQmoIha2YnMR2ySuG3Y5WcTsys+l+17J0
nOGGYXYt+HtZTPCVb9YW1ecgka/TygoZnSZETxTsCTdaU2BMkUTMMLeBE012/d8l
oQqt4shRjWlLi3aVbEqtjMPzFJJpAYS3I6mfSr8W/LQwRz50NGeq8fWWS9cNjj9R
UqbztIFdZ26c8x/0HLAAngwc1fPv0gDWfLDsprJzPGCGb9KsLEpRJ6JAC4JY8PsG
ndq9kcHpaFnVxudo+/XmUaVUrEKPtvCaDqKNaHZYlQbX63O016l55Pl7pOJMFX7c
L1F6GJOazsKSbKQUOXB7BEsKtcQi6InSycFXc91Lb82e0Cxx1rhxQj7GqjRcD6ju
bPII40Q/OxLM4N6HfEAM/9QxWZb/GUqG6gMDQIY6ygXP0QpLTWHi1pj9F/40o3oa
EGUjp2fpNDhWoMWUtJumMhtSnuCnSXNM59ailaqcvKDRYa7Zo+yoxmGiu0PCVPoN
W+0+/mlQkbG6Z7vkta0IhJvmzeB3MA6LixjY3qE/PByXrX1rYc6qAj+yRWUvRKey
jhJf/W+9e4HgfQ31LEf6r35DvBPyhySlM6cjD6Kr5/Q8FCR5gAM4QPOt1kOoCIJP
4Fa9YpXrYcFRKacjsbqHVE0owWQhjLLKIAEK+NrOw/udNEylbaM7hVpBo7wdSrqd
QSNJ/LisLt/zKPCoWOU9LuMZIfrZwYaFgzFXnovgdCCLx3EvWUk36fMb/YAdF0Zb
DAHozSASyejh7LBEszfYstAohnZyVV5o/NJoTif3Pm3JQ1xi4R+Hzhvco1Np4ZOX
v9vf//LKMVkqZKFxq4DQhCSaIF3whHaknxYbuHTNy2gPZdQLZHjWa1ELNuelq1ks
jGvpFPAY8IUg2JSV6SWtnMTlBXbaTsZL9YFCrbz2mlqthYQyZbxVsZUleHJT2LN8
Hg2taE4o4us3ZbBLU3+RcKU8lMr6mkDzQACGeAsfJjx2TdoDBedXOn2wPHl/iMiR
jDLSsBX54/NYbIhSWJkqjbfhIEHlteJSqLx3BHJUKTNrF3SLRZswICCw/2wtUWr5
9AUOMJF63F0XXNzwC8VP5N3TWDuO1gL3IxMLFVGnln1tyEGuN7xci70NWlLbWTt9
W1fcjnL56Nd+BQgCh/RaoELQi+Q4Ju8gvtho6/fRsTs8K/zsSEt6k77zSCDCNswR
Ls6pEEdjYH//3f7DwwLEHWZZj8ggmH3DP6T7FclMa0blGFN02+Yrr0ki+NN+r9yR
/bHqIShTV7u4QlOpK0B9QwLbHr4AShmHweKX0OMgL00XMy50rNQkquXYXa4ej12E
5xNabivWwYQtS468K0IwNOtOd3+dZ72xQDFn5N56sXklEy5JSKqejx5Em2r+3sbC
RISlD//+VlNbw3qmq7I1dxGRKB58KkogcT4DOw2qDqpqM7ZHGor1BTbehbItxeOJ
03DcNrLyDQMwSJ486WYzYP9gG0f9tloVWONV5Tqps+mr72ADBKRRRSSnOQD+XgZR
+E+EBPnK4Hsm4aeT9MOucwj7ymp61EDXd4HaVcJBSrQRr8R2ja2gbkWCi8HXbJcZ
8odvhdsblaTxt3SDqSJlnY0fSq2XIIlDzrArDeWgT6Kv4DeGIMSS5aT0+s6UpNhI
cae9P6oofQ/2yRP3iVfEXOGCXLF9LyneELe9uZkvgoV2U8HyzBheoPLWzyaUgLDC
bjETyu1HTfATHovTU0ZUOptINAN/t8WAyQdqYYjXWIqWfNQBYLSoNGz1Y+11CoNv
qSpVCP1j+3LvxCpuekpQqeisKX0af9Cw1FhK/owCippgUaiZx8bKzxnJq4POAYjh
JOBxj17/YEMlz9EmuQ2S9o8a6oSv1H/Z3n+YzCilecE7DT52/UF8rGBcKBv6pqbf
pHV05Uxm/NTEZ30P4g9xEvmaDM8Jdt+JarFpEWNARfyopTR5SK2bCblgAXkIW/0K
a29/NURS7yMMo5mX/fnWZR/CafDtDG6d8jt1llWSQoPfkDH/9R60rhG6byz6xeYe
NuRNMBsWqr8bpavL1IsBs8P9O23NgcWVsfBxVbebJmHEpUPvEqxw9oQNoEkgzOuq
244AlSd8mpkb6UGStFGEaHavE1H9fe1qovHBRboRHwX9vTOnYNCOnUIH+TQo1LzZ
bZGDQOeQogadbHIGuPh2I8yYwVDpL25BvdK1wtqyGtSYocsomEmb+8QQoos2FKcs
ktYCD2yO5ACZ3Gxwk7mm/L0FUp59DfOpiyt4ZwclsnPBJkwPB/b3TNya+CrdKc9Z
NqUtFt0ZOG1EXB6eotRrYAuNbAv8lFmQfn0WeKDUJafoNtPnq/pSkmc4GS+h8zqp
+BKoBS49RNPIhKExvs9OGN2v215eAtz36ktjGYBLYjHCmtKaWe3gH+hfxlWIIwkq
5p1nAIesKza2Ck+MTnsq7vmPpia45QeNLTcwsYz140DBnP63VNEOpd+5996T/c9g
YOvpUdyrHnpP3SrX4xjVZQBnqdw9/+1fKEUNp413ahyLlETYsuOJX4Bmcx7ljV1E
nY4hxp5nyVjXIjPSug6GyZkdDe6LarBzSnivkHkI7fuadR7H/PSUQ46eK4OzBE+i
xcxwFyH42vmtjnLPuxIw+b+O1ixtAe1jnklW5ELC3euBfaJNYdu+Pgf+0SyUPjhw
2E8JKHKUc/KRx4NJi2eb+R9wH24LCVbzC1vL6Bi89g4BpT680Ir5cp+aVNDMsSJb
x/KhSGB2b7QJT3m42br+LvFpNYXzb9n7riVsxgnBd0rGoM8kIXSJRKtRscZQ/9Lc
pRp0PI7tXIkHPrk5RMy2iQeE/Ek/UebqoD6D6IlrdvhA7qRRHmrhcnEkaTrSwR9V
NAJC9WERENLteqFaevd8gNqxU/kAMhij+xxpvjnky4jXmng1Pgmj15B+1yqAQwXu
Wv7M6Zc1Z8BhLRrohxPaXeZ1b2thXqR/8kGkk9r5/KP3S+fp4P+mn02/+0kgBuG9
1gjIz3WtoUZuTT/2IgsTRPSu6T+asUsQ+ozEylzip1VafuhHTpiFgtXpr9qgO3Am
kE5DyuJUfodVZ9Rki8fJgImgVOBnhcv95AafnkP/m0C6jg+qnXKn/+p2WsBldVQi
itQVp/5R7zI4hGQRFyoc3ail2yqQWfYpnHd35XhY4Kl3shQUqGJ5UJxfUBgPkdLS
riU+/dHbkyTGq5/4/dyt/CBECpCFzA4oeVz6bv2YNaA2woKd6eQhx8NSy12NnoAQ
fynCz2vbYtLoY8QBa1FYxJ1M4Xkd5xB7idPeqzxPOggceLCD5Y0OB1q34NnMyCxU
a6YufKrVr07ooWqjS91DybFQY5i+UMeS97jnE0ILfVfWiw0fFnTF2nYU2mvcGtcZ
/LJNXR29MgM0o5PV7lJCPWYM+9IPkaR7Eg7+++zPt8SEr3zUC2Qr3RwVqcpkxIxq
R/KA5mbddQMPllXY5vcSa5Ugd2gFGQroFkU3gs37rpVA1tME8MRBKjIgA2yzQ0tP
F4+8hsTlQxYhpMJOcW3rkSCy13BHnLh063nRQJsbdf4mKwJaTrhQ/zkw2fuUr/vA
vjUDTdBNwyb2vm3xR6H3y/Zo5jxpSPY3sMaXj3E3XqKhMIh9JYK1TSzMFhFDy8Av
zRvHkrMF0oIyVarEZLyQuP3gAYkXjcfOgwau65VehLgxULOUjs8iuNXlfp2EViT8
Up10irVKYj541HxGgSOmjA31NF8t4bbTt0L0SZXcMh69NOImkwJxpKK84iLL/wOO
9AxOnh0IxK9b8R3/B7ZsQPCu8n+A6UtSKt6aQ0v7G4CVQuxYPPDWZikoha1Hy69v
7Gkc+3/PDvVIZspcHNm6zNjfW6sjjhjY82KBS3YkeKVGDYnaAZd3h1THeRvR01Az
W6ZHVJQlex4qLw5c8l2+HX6BZpGfxF2ng58ONZkcAirnUqLNu13sHQJkcf1U6c43
TQ5PWCUTEuQ+hoHOL9YAZM9NZHS4F0X3BsH5+qL1XSWLfYC1C0HsEgaQX+Ee+M2C
rJwM//B5xjRYu8yH2tZZT9O9ST8/mpvd69ffmkd9dyaj3aqXZ5vJGp7t947JeJod
ADW1J55miX6zhO7BbdNvK49YCyqqT0WKsIPJ+KQ2iYzlws3+XjRvuDro7CElfBQA
fTM6ajC44/DnnXUjTizZyvwfchseVD1YnCNOLgI8X7MRgRxspnPgLPMuIIpebqGX
YSjlTqQIN8uINokppYA264lJ+bnc3sI8wILCH/G+FaOgh3WjPNsDpGnNsTDSy6oc
kcapFgmNhOYSPt4yPDRpqxpFM5gJlujY/a2ST+xF2ZmLPQKJv5lXCflS6mRVtP1S
JR1z0UH9cyMMnq8gbJpeyPVMj01uvjK3WTHnzKzxZen/e4FO8ZFzqLrtNXw7ySyc
+0ofzXCvYr0iNe+8KH/5uKqBbTHIVMfmGDgLNodG35ey4F1YvZ9e6hSBPaSrmhut
qHWtqlsPj4frkL4k/wWCg5akUvfCYgBx7yIFiqmsuQ2D9ceYo6cZ8o+a/GrSY3P8
F+AkCi52L6Kmgyqkp5UZrpu2lfQiB53o/lNQHLAfhJktEMtc2mkLSu9PTApLwxd0
kQBE3GINxHyZTl5iiAKXJw+T/MxBQRKO/q+uZgKtxzYiQsgCQhe2wn55rwQwF9by
hMMxUC5pDMpQl4e58CN47yZJJVulNwKi+DDf0Mih1gZpCsUcNDNVC9vVXXRNOKOe
7fHDvgvqNC0ihjE9yVaJOT4AQN9Msjg9zJSM0RT8O2O+1x8bWQMQwKXgbyYtj0+2
GTVoGIWShisWZkA0KUycKgxTVtNWBn0o604Dd5PJKNsySOzekN3Erhoh2U+vowxd
oWmmKeRF2dalLDpIOKOEiuhKUbFvEPV6YDurb3ejmVX6ahQYZ/O9tqK9GPwfHLAg
pZPwJWPL3Dt72fzeXwmR3Yt7WmN86FA49sB1mpSI3ISr4W3ntFKeRPdFZUc5Gj8w
I4Davqy5MwWZhX1tPIbuST1R2XuFyqjc1MbNB6ihwyygVCPQonZ9Zfe30+jCfig3
wgSfqwzfJkT5pbwUROCBgQGlS/iNkW4zhYUfR6RL0qc8k2xpaaCR1F4Xl/R/Skml
doQd5Sj+0gzHqAr3xwKIz+pZqcThL2IPFBU2YQWC1O3OVK++yIeqXCoH5rvMySk+
Lw9nm0Ah+1+fKaeGqwOAggbvsB4SP8dOPh1Qo0TkimdBKBdn6vcxAlQWq87ocsca
xrcwcBvseaO2r4lSX+zXpf3byr4DoKqz1oatlD3KIMDRdTCdvV0qaOLCDIHLwKeB
Y5TFbJiFf5YluXKuWmC28xJKxipqB4zHFVrfcmSOCRR0lzzMepcejHoD5BjBPDrS
D6Zs19KQDS6Q/C7JdHLQH43Rs2EuJ5e4Vy44HywxrNYhO12d1l6fiFasmvPR7snr
tTj17HIm7gY1Bk9C0wOK3k7tmSLhondVWwkDwY08S8L0YrqjT7qDXXyESUxNBvT3
rKFqWVOGI1BV/GrTt5+bR5nz54edcxlPTKtN6jTjPHBiMurHLFY0J7No0cJOly7p
daUr+M7PrrsZJ0uFhlX0qIYtRMGu6MM44eUq+0VHrfbVvAmfRW/JdYjM6u9Nt3ig
wpk9P3MP+h11pucCGvH9jVs07Am0SCRUkg+qJznQ5i0kSpefOUY0fxGA+YLP7vYg
javH9sg8LIy/p1E79pnJk8oRcB6ralsFrCSjHU97S7TDu54isLRXH1ueBNN7FnYJ
wlFj3Jq2Fwx6c8hPwij1KU7KDeU4394wvBl34x8VvAovp95Vn3HOblGdavgNQoxV
PicA/AT4xMWqcfhPiF+gg6eU+lp3jD4wxPptP78urXuhUEszJyaddsVX5FKJ15AM
DJsjBeUaIfr0IscRXtr4dXSPfnZ6qm9R8p5CHHoerNLNtWdg/1XrTXWRVPNY2L/P
/dheDJOeGMk107ft6SK2S8U3usgmO8Al96UysiE2OR4BgYp12eNj01rI42GrswDq
YE3BJuNu01YrcYNCcPLW5OVILHPYP7xClNBPP21BcchRuQTa2zti/Y+NwgVSGDwU
FPkkZBD0LsKkrSLxAoP7Pkfnph5LKZ78McVJFxkNHKNlK+KOM+jp6AfF0usqZ7Te
x4HGfpbP4PFdObQZXYgKYvXsnb2E30cLWqCSYKTSQv8RRUg+QSuOVnka2DtY4Svr
sMkc6590GyQDE93va2U70HRZUsNiUrdyGA0jA0TzzGbeFxSnwSc41az0bK6J32fw
Nq6DIjvJO37eDOyB9FSEGbBO2z9utgVCrdwt9QJ1+XwJhh0hm4/oWEbD9C/36JLy
njRnuK32CFrJ4zIPkUy3F4yd8udsLtPIF9Rztpn3964+UTujeX5csUX95P+pRXba
IVaGeal2L4g2RzCXmYdAoTHaDszMvgrwpMb+8xLjOOT/Ri1yNXRNZsXIdN70EUBC
z134VNZ1gKYmUF3HKWzQHxr71O5bvpeyD3RxMSM+WZdrViSHlkowynZvdOHYBl2y
/yoP21vvaEs9qzQXdXuiAjtoR3Yr8Bwc8H9fmNsd4/fdGcwCKDWGLyDV8daNK3Lm
eofqR/EjzPZAm4jwCFxPoeOGJ78OD4BLszhetp6lTw3xQjNaD/t3Ns2IiUBDRsdP
n07dFIeWEibJW43lXRbxUQwu4JJ+X60NDbPfLS8nyswCrY+e25+FordaAJ9rC/Wd
EP49EVHc3WAQO5ptt9hRdQiEhGOCq4t8kXwz837Z5UHVhlzR1X+eVeheaWLIFwhu
RKGtkyn6yLEOifdMMF0EK/pFiNESDGsFcQdIselbhhR4g8jxH20D+W6gnmSmJUWu
UAHXIMOtIDyyogPDiQVVAqssn9wt6gm8FN7jFbQH+1SOMZU93h6K/CuXAqY1YrZz
mtJ6v8ft4QvFXRSftaKehCNd4/DiVSWLuhtQYRrVdnpHsCo+nPmFEpo4rU7EgQLP
mK8aAWhZ6cOURFkdi2HYfJv7UbFPjCk5RNn1oiEqo/8AQMokUeCUkwB/xoGiAMID
vInZJZubPkPmpg5bS4megoT+ajtPGn0nWShGhRMxHV2mNKvGdIEiyrbJhGp/GCTF
2Dttm7QyH0RLAlozDFtVy0Gkrku7yUaOKkFEo0bdtyxRyhG2Aukeh1pGcNu45Ya4
7XhAZ0/4AqnMWZT0Oq13DFTUkyzIdGdBj5fBX7Lw1PJc5Ewl3+nqeK0pxopx9eqa
2Xz0lxNi82zzUcEoJ9Jt7ERtjjvaYuEcUEiDd0z18DByKRiUUcZO4PQgSfEeD7tI
4nfZa/W51rD6JgJhakBK8EwGWkzWlwIq2CStOq9f7fKdY0RcyaFVs9Qci0Snnq8s
XNja+zQYK4V2ji8VVPWsMCC+in9btUCP0DuO0mREOJuonSYi7b/ysI8bgKLExmF3
xMYCFrQmNI9tGGDaeiqTj1MFPjGbPzum3U8GSVug6XJ83ACRBweiisZyKrUklxtG
MVklIrHVpTWN8Rgn4Nb8WLKpct4slduZXrnE+f62LNpDiOV7k/ElaYf71RioNlvA
8gSFUCkBoIyw6zbfRIDoaOd58QZo9PVlRAANzE9cgZOKUUbcUN+ozzo1jZWF2PQH
5OAgubvyP/MEur4CB9Dig3EoQocZLde12SmMv84CyXmvjhmVMkmsScbMrLPVCHEs
wLHptsfl0bmlPzySIkET1qvqx4mmSKlIfGyOTcXI2lktKBzZ5pIKvitXt16B8IRX
+K3/vIwIfEtQZdLLp5smSknniQ79lrOQNjPMhRzxZ3KyQkr3V6jD09lENu6iXSZE
xX5Dmnz2XIaZF5NuZFD7Yuput63WRAMGmwvHlRFk4FC/wqYU3I9cXx9dRYg8Lapl
x/0SHMU4eMk2D2MtOohkAw45Wvjzpw0jBoIXG6b9LP+IKsZJwom4YB+7oTbw8Qw2
Mj8SdVAm93qiYdo+ZqLUI/gVo64d7kBLdwFRZ4sPwgCwJ76Hl15S6NSFQQIjZidL
tVeo2QNlXPJPZc/3a9v/PDy1uRCRkdAOU3u+8mBJcPToEB+9sHaJe3Aruj7b1TEo
Q7BC++wlNUDjVamSKwMUdhjZZSnl+He6Hs3yYxdqODP6OZs1SP2fguxsKjO5SbZh
krCtyWxmv+Z9BU33q6BDloWZMSBabikprg5WLAZN5JyRsqSlUSqXD0mY/x/fsGcf
j3ddXJFFJCf3XYOwVJsZJX5d4QVSIpHf0cXS6D7YmO5B1EoYwHLCxJgBD8wEY6K/
EgBbDQYpYAvZQAipBpfKnRrx/qOvNurGyUPthH35ygPNmyCC2NqHSjKw7+KoDxjb
9tu9P1fmW4w8UlWID6FZPIYq7Ab8UJerkhSmtpUI+4J5oUHSoQi3gsrx6xUcsplh
U9iTkBMnDWO66XveTSBTfzVXj6h+0g9Tyb7kYA4ZmNTAxLCAE2T4fCA8eYFgWBV0
Zk+4duYbmbtWXpfmPtQBjdjX3Q6FFWgsdEW7Am6QNJKbBBxXyBrsBYa0Bx3eMfKX
p9oAJICSdo4C6i8VdiAh5JJc5uxdyvqm1cDi0QAJnP54zBbQj4oGAvvmylstor4l
o9eQ73lMa13cUaei4uzT9zT4QI4pQbGHCTef/+df/V4ZLJqSW2H+XWDs8cutVsdp
qo6dpUmYO5SsEcMSRCn+Z0s1J9uJ+qTWiV/QGueSOOQYcSGeOWtY0mF1aC+7N0Ux
mIMlaVe5ziGX0BqhhNGeETLSDXhzCKSNEcQNRkuAOSCMLmjLfxkZHqnAhpd06Lvw
T5dDf0iDqyCv+V8x12oyZpQAgDlW1/SLIalTWLiM4eJMZjrDXw6kn90vvCU93uiO
E6UvxhReLAPWKE+9CbADut0+FgeaQqfcm6K/BbR6DtTuldNGOhKvPVXMwz71gh+a
LbhnvB3g6lfjZha3aLcFtIgipZKOrSzgSnS8RaL1QC7UObzLueNbxxtswOcmTL/4
vc5aQks+nSXAPfYaz02evJHumYMqvAW/LyKfXJT5WIoe7WTnR7lJtvi0S2OY0Oqq
pxxx4OjuYTfAKabJsHSq0PqCiRktYX8ibvXmxjLZnhT0b84qInHXUUiznNB7NV0o
E2Mfj2ozQ/CTVewoBUi7zwIMbEd1MgkuPEZjzMXuHQddiJm1La/D6XX2G1AH+6Ht
ppZ4HHKX86J7j8dmqjfIL11OnWXOKCY5WF3+vXoCTeYQ0ckgrDi8+FoNKYEfkpXy
/qguUPvyUT9p6DUy44E3loLYaicjS8+M/AQuPI1i2OoB1m5T9S7X2AH0Xfq6il77
BFU4txn6Fz2z/j2pkkyhISbCNvzUxFhFAB9MNV67UhJldMWRPozp4LMjcrQx9sL6
4zUAyhHDiyRXdb9iX9UaLNzgzQIC0kw2+ADOGiwBgx3YgVxUvP1h4ZVAlhGJUrOp
sELzitZXiMwgM7a0uPqvlw9kFQVLVXm6S1wToBO7rwlcXBbwKlnfIsXXof74j5x6
7XhzQRW6VGjjGCZg0+IOVJnLvV0QGiqA4wbD6zjSGTRZxFdr+ZQSaA8Gh+zFFQIC
hPEtgsHunoJq4HjzBep4Gs7gaPND5awpnrpxtJJ8kzF8yme5AR+ssXKRCubS3TjR
zAcFA4Yofw+hZpQa/Cxe9JIZUatpA8yZSA8Hk85LLEsFXbSWyU+J7/nKhIipglP8
gTXeq49wxiKgjo+YBxUW31qsyQ8FoCr03Nw/0lZICaa0DBXajwY8T2VmEIIzZXhy
ZvXnRpoJbQfc39O8ENQxZdMknk1/YYD1kaVKAMPF5DXrHIi3kr7xoaDuO1em7z3w
JDAyN5fbzuSAX8zpGW117bafKiv23C1pwrBXeSYyn7o6A0ouMAgQ4aDZ932MONTX
UayblRSd9crGPm5fFYWpaD1r3oDI1rYrj4gxzCG8l6/1dWpoWIP3nZOhcKouYMFL
SBaM6A0oxxfJKZCmipNObLiQYwsBA+QRhBG7NgS08Sbwvj0OVDcTPy5YZcTDX3ux
AaEwW77K9N0WfeelHZ3Kw8o2CSMrLg/SJsrJSAIDEv3tYYBeKzXcsFZJ7Wjj1A49
f2bvNFzb2eA8+TtfQB8Z3QRGGjbaGKgz2/guerBy0qPBSVGbczK3244uErQYCX5V
nUCTbjOyJp5xnhB2Y38PiN5XZnEMoWQpsJ/MW+BRp9Yc4C8D8n90fEWB9FmCDP42
RsN8KzrZfZm9gcgVgmHfvQobCp4o4lGWs338NBlTLe1n59HCfBsA3Bcbhnflxih3
IE1Hkwm5IBaFHaJwdwuGx6mj7wgL5a9y4Wp0aJw0Ey/VNygHFjKQyybE6hR2zqcz
1N5IBAnbAqO47y4UQTHuqX0SZSZ1mkn814Spk0KSD6DH3egE3NpwsipW86Ff6XWP
N8fjdHPpIFyv922Mwh3k4iL7GmK1xGqiJ4LICNN0n9FcZdRBNeF5VUMib7QAZMzu
eoHyvRKzbhMpd960VKr7O95d+O1mRnRhWAyk7YfsWITN5QBB2OCuqU8aTqTFpdG3
w5rvAljnywbewlqaI+z+u42In4ttu/cALHqSUKCixV4JjwSYeQBl0P3KgKhfc0FN
d6LazoNVcHmQE3yJS5GblWAYWYBKaZg/MKaLP1uTqlKV76gat/0aV01WeXgJhEgp
L7v5NzDug9sMOmvI+N2z1npBCDyXqT27tBo0PSyJdf9eacWoXAZ5gOTzuyqHaJuu
b3Td4+yaDYHx68WaicykRZzFvj/SGhNj1HhU8o9kNQIArZlY0OZbCErvk4kbrjjq
wdYY9xqLgHR8VKfWUTMpirSRNgy+DumgO3k/xcWpDuKz6igXZC4K4NZnfDHpmpc1
fn1jJpe3QSOtDN6jURPwsctkJ2ivEisXblsippIDCul3immB3JWuwwAhasmMqGzL
YPhnVby/BV1GcOGRkPrp43lCemJZCk67LOr1SE6WVVSY38bWhEmgIbU8voMwFZBD
c0/0PCdzxH2xeNdx0Rj8l7Rx016M6U6TRCZy+2ENpvAbSySPNRV4SOO3XEQ1nAyt
a9HXju+XL38pQuBNqC61IwgH7QRxk3zr92aZl7/D0VV+t18N6rg2dgJmApFpjxlH
XBn7kRhrhftvnibzPiZXNu8faQ6ksNimIKtvIFHmSzniWr0rjX7Max75tVLf64AL
N0CqTKSnjM3/Gp6FeJwlc5zYxOam+2HugE/YFiRjkDpxCEPr1Rb1RKnaj9M9yBKF
9CZmCgF2lRwYXE3XmuT2GNeiPcaXcnzwphByHlnJbJ68hgq90hPq6G5i+hsp8NqL
zvjSZJLYgX50v8AqdGDxcIFqbmJUkqyPUs8wSd/2WkWc0pQIV7qvYAEWhDNqk7dZ
iTUpSJ/4+kgVg5r/EQwEhBgE9lCtvIAeYjFcKOEk9fFBoETx4GEWrbrC9Gnb7fWd
X5pKyJWjUXplzx3LkJnmpqDoh+deAfI4r7S3bvDXuogGdHX4Et3e4SNPIvzHNrUz
OqEkp7tfjAh7+QxYa/bWabx9P2XZCHYS1AsyfIHF/o/u0IOA0xAZldS30OI6lkNm
TwNcKwxUjTahNWGeFmT2ldD591JMnYBfQwqaEYjg3roV5VYqMD0/Jmjt8VIQxy9F
05Cx97hEvvMp9zwm/CD4aUdtm+XRAOjweub3zgD7/CkCRVvTFDY/IquhU+ljsq95
/5+L/28G5kOamjrOSnUmEnp0fMX2dgwh6GrULe35Trrww6o+HrJF93oa7aXTxFN9
WlVJBqsFtakMWQMINqvakF/ywOeDKk8CvWzoEIL3/wzN8PZpj8xw+4IHI50GL3Jj
3JXM0dM0fDGvoKJyS3gWBxhVhhGjAcwACeFm1Lz3ku2+qGltPktzm17zmZpnbDtB
c6via/AeaWV62PHn3vyMlcbj0nRnn4SPSra1F9HSMJ9ECY0XbEnd73//3tbAbxIy
skGm3y6aPZVkoFOb0eN/GWJwiefHmUuDoqMC+UO+JCYpapsn4HtKi9G5YsjzwamG
pbPPBv0tYpLuMK7qRVIx9wKbgqYuchGqyOmrwOafx9pJfQzJQhaT+P5XS0xkrDbz
oX92xQYmVudKwa4C7EM7VpMeCuTDc5yaNLwqlHFH7sSqcKFZG2vx7hHLdw8uoEj+
tXDtkZvFOEPHUskdisvOTv8cSVwU2Z8uDGM3/lwYuFBLavAiwEiSUyDkiZ67e8wq
btntiVLa6cqDg5DYYy7bPba/KfbiSb+SIBhIs1vMlOfX1CpXjdHYB6ONT4ZMZv/k
C6pmM4w5dn7Oene4Hy3bzkp6bWOq6PmdydqHcA7gZdhWrfSh1FVB9++oMcFhIZ80
fLpX3Bf02vURE5EaU5S7zkRcWxJki+ILjko2WOBivCcT5Yru69fZO/nuoue+txeX
LpKjMeCbP4/wsuxMWdRxdnL9kWCkjc+leqhy41t45JfsZVb+ludZPWOehKKLTndr
Yjp2/UrlgdGuY5QEfts9ZL80gZYqgj9SeBM2L3/+v9jzjbmtA0HQAe3oPOEytzH2
m1kkT5qWIiCSwDMW7UZOoGwxfEsz/bgGZFBhcpzp8/2N+nM7AQ779vjccvI6nZXB
V3Mdf3P49O3m1sd7ZbRDlRdLlw+Shn0QvWuDLv4WivZ/90C/51hHWSSyEoc631BK
2pojq40naehjd71c8wdmQbbVVLzA/icWK6HkmbeuCYD+qQ1DlM6sVueWAyHBhB3C
gG9DALeZaKiNj2sWifvZU6Z5H1AGAaEf+UVjBig3hWsVz5nLhQnXSjx35ufV72+0
OukqmeRd0uX/z0oDfPqTAl7su1FEvHpxHgoa2mQqVXJBxHhC0xM+9jQbSR1r1gUc
Wk3LPMrYTvriAqXi4I8CmMgQCR3N4DXlLMFwZIW52iqi8JQyQrpT4hxlk+oMSYzd
HM83lG3qabOYLNMzdMaNJUhRywdL2sgn11Y0BNB8a7UxfyBRWo8GSyVocjTWNlro
D5aMrLxdNczaGNa8VwARto4HkhqybkdRV8WctDkO3SPlNos9A1qJnf5rzxf5sUnD
fsfWs18T4pXlB8yHxrNW/gzLH8tZ8wI0Y4qWrlQuXw6Cy83W3jOaUMDHyHr7ZzHJ
awtZPaKeABADHfEyXCBfM76QNv3kVQdmdh5iJQyBTXxJmHBS8SI9+LCQugj22mFD
tlH8g8M3a9Nutp4zBj251tFegfJk3HOEGwjQoavuMfXEKLGx1j4/53jOfEVeAUXZ
ps37A2OiNqEmvEZBi8jkvSKRWcU2H8EnIKydZVn47mqntlQ9zM8kmKUYXcqe0V0g
8bzmdYqV5ZM1fAg6hTq5Y39Yom6OICQG/65f7uZXNBxp2/uBd2ly7khtZq32rirS
vPxp7Jdwf4lyKfMV53XKzEDBDHhz+5bBbTVSmxY/GIhPBnIJr1IeQ0gCsNT/GqD1
JPIo6stAbaqAwv4EYe5FzQ4KuwSSQV5lmvpDqfb5VlbGBVesJkKuFMaMOk7IPXkr
mtkH/z+9EUjcESqhs1A/mqot1b3ex/puob/wYN7CRKnAwRR7WAnaFBY+Vu1La0zd
xvLTO7P4u3sOQq9G+ZrAqmSh0mRTxpsNixjYjKdggcfQlHFfyUgBZZpO53bM8Joo
yqZsKi51dT5Y0QzcuJe2ZHoiwOnULAzypQRKocIGVw6h8vRB0dk/6FzXliVTruof
b/pvQh9nsgw/xr7SjV3KliBi5Tzh5CHo2gXxpua09apo4kMfwXjMpc50/wHpNAZu
7clzq6jCvjLS00AQbuZlYDhb1oxYbTIXB8vNLiuqhYmUwB6vUaYEwQ8e4w9Knjko
sB8MJ0Ec2kUJfSSxraWdei9/CYm225zkRLiqtfz/qz0JQOs0uGjdn5dwON6ho7t1
NCZJHqSDDKG8JNdwNRHkr8DNNcTMGJpT2fR8K5/I0AX99FKYYL8+hLIhd9sBMjou
jgybEiZnDGX3ZF0dyJJFP9wlK07+Dfm9NZIw+ur4pJCoWD9h91Kj2WMno+YphBjp
b5vTzZSlAhFGPYC5Pnuvg95Kpqj/tNqRrcqY1cidKVXkq6QWbKTFndzUdCk+jPoN
7i5UPD9oElr1n4qIJ6B7BzKisL9KFYi9yiwCp3Udp319JjgWzU8NAmWyx8AZd5zA
e+e5nvEIxtL1LQxNMFVRehdrH7OMXExzZwSbtJP/K6W1hbyNeNJj+vpyu6yrqFMQ
3UIvZC16FG9grYZYB2j7u4jbtOK8nPKVD0rotaa8wNzGmqzaq7U5z6mUfuRLDy1+
quQkn2dVydb+gAFPAi5RU9A4WtO60DznQ/z3uJN9N69+xpGE7rqrUBiBSRRzRZsq
gaI2iQzk7IqwMkqSO9NDrViqFQeqFEt5jValA16YHXlh8mejdfNUvq9JdDNMYl6K
itinySw5pc9vgPxHizcF+yyUHllMkFLFBAdJN2QbtVJ7Jx1y+iAVWcNA8iOR+4Gj
mJxOXWoSL31Eph7qT4VfMq0R79ieTMHhrH6y1tAAOVvGWWGS+3FaDwWjTU6OjFgx
9LS+T1UGOiN+zpvOMlYrAgN6f5fqRERn/RBJM80pS1UUrtso/eRVXqRFt3ip4QF1
LtThomiXfP8RUFrld3dpdjt5yscMx1atlHMqzbyPxO2YGUavOeVJZJ3QulyqHjDs
bij31s6EYFjd/8TRvwSXSuWzGWNIXB/NLlWzbDWgkcjlJKFQLTn/s/NImSazb06g
r/T7aoS13hgd74pWYaaAcxilW+im25Zj/VJGkoJc3tjcYdcprMkl87b/gaYvOmcg
KkDqxeEKXNDQJSZ2bcPe1cBXvJoivjYBRYCsDlKZlFvhN4lnqeCebASn4GvwgxGG
VRA5s22WIe+9ec/+Gqqa3xP2wGdUTLa1+s0cETTEzma9xVxWq1epwYKC1MdSoJFc
4OtEvA7Km6gqZ2e4UcPvMR/nObN2FbU3GFft5nu2S0GgTqE5HaR0ogrnXluNyWNs
KL9yBs9iViikPF9IeViaT5/s4o2Q5m3gPuwh8tsYA8DymI/yTgQQHRhkmWv7SKjS
MCixBOCpodalXLH6Y9y3/63nxBjfHvgMdvQFLNPLwnlShDgbaMg2DACe6P0+fiQR
QvUzS3tr8t+NRB3iTd92ubWggaGBqvT5+ejbsUC9Ns+NSfM9B12xmKQ93W+Q6aUO
FQEAzs0D9Phmg3e04MwPeuKtPt+o4lIK6g3QgDgdrgMTAtWW8dV7caJrhD/mKpVZ
qhK/1xDPAOp5eBqg1g0cqDrGP8HvHenctE+XBWfAT15muG4ZRILrtJ2mSk2TYlzw
NC1y7uAgClnbehp5nK1KWpDSXRjrMzWEXbaILsRkIzlPgzeaFhmqPF4BBgznmr0i
99kdcbpsANWvhbQ1kdde7bQZjVAXIMwUIgGcrbQhnqcqUHHkA3Dm8AHZd2+n4dRV
CFZMlko944ULcMIezJ+T0r0hjcr/FgnwFVRaNsdIFoj5pCM/qCbOpBoap9dmNGrc
GPluqwrisI9NP6YAu4/zM02gVbIpVPPFkz7aDZdLGOfpbeLdBVFgHMbl0KGI58NY
U+M+pql5P6ZCgs3KU5cCcRN9fna2amwQxVV7FyyPex2X/ycDbntTNkAVT84r0sfj
R3iJAcD4Rl2ER2WIfCEH1m4P/+DAHSt0YJbHHvlB19S2neoSCervjFrj+cXrk0mi
BI13okUPwipYlKkd/hJbd5rfhRcc6MEijtXolUb/4g+hoM7IwEYebMulRw7vikh8
Bp97Xuzus9fhjvutkJF/RCfhpZ09ZX6kIwdvstmlXtCloxDu3usIOZ1BM6/aXzxR
JRt8IC/X4HfgRjsNt8qPC1VzgNOtbwKBkdcXrHyQHvierwfrafOmoe59RMepANAv
553DojS++dwls+zb3pu6k51SIYgYt+J4mwH8H5AlUYgDxKnaWh+IeI1JyDd+DwDx
9DKyaDXd8e/yvsUXKu4JY42fnUkS/5oQAI5Y6Ft1YNscNPgr0/km331N125gMhLk
t1wOIpeSsm2eoAlzmUtpDOX+gXNuLKqsU6CWp2sCIuE0fa3r5+WyU9hZMH7oOemI
l8cg8V8QQCHJLbpq8JsveQGwOXeSAfBqVBzO7qV+qC4gXXRyll5zr+ypZWNahO8p
RP2n9OxmArSn76CpdLFQbSrlX+GdqRuxzLKB6YqTrJuv3HBroEUc6S1WllZ1FQ3F
TFD7EGd85A4j39F3LNHNaPauKZYl+rOB1JvA7qnDQiu2VNb0bKd+JR027yVkqaUD
r7mkolwFADQlexYmKLN92BcM7hEFq/ouSfvhVy6cy+q13p7MvW7tn0/Myao0HFGQ
pqIZmwo7D+TV4moVFhsC3PxYpCAdmDXZA/SuKQMGECldSgPDkajKcXB0xtsIVrEw
+9udjlNIu2AcRcSMW60Zow1mUzO0lAkg0aspdjvP+SpUUP/f4AIiMvj26r/H+suI
ZqTY4SKB2+qeIgqhD4/ofi3blwZYOrOa3WyPjr+4o1yrgfEbuXBD8yx9jtDNDMAt
AcEpqB3uF+jjUMy3pW/mpdEQr7USyKJQlCkuSGTZiXUxxnIoNGv8byepCYMCIo1M
nJZi53pUp5RMmRDNq7gOWB4fNJV8PA92EkHSstRi8ewleorOkwSe5VORXhDAnwWy
K88j/7WhFXIb+XKjnVcMCud4HZh1ikjP98tO4sgAfPIpFZ+elQ4Z1KOJwHbseKpr
v/zE4ITvoqP7QiSfZQmqd/V2TPH1Oh/zjSgmyXHLWzY6LCQzU6nIJlbmwwYoWDNe
/f/RPpzv2ZXuKYlmv198fkc5aB061OMYWBA+EXGhV9U8ViOEsfe9VCBUn9nC+KRV
Aw3taQQeYO/vckk2A9VNfSYv8UCZy8D9RVZmBace4jEz8B+8Z881Q9ZTzN6pPdct
RDIMiKwgGnBqZlT+1ordsWweYYIkWGMtWaPIidjbV9p2hPS5GlZychjCnlO10x/w
HUp88d27WI2LLMMrMCtJtrAl9yofPWIWP1yZoqEfbnWxOMMBUAFX+gvzzbp4Fd+n
A7WwPhcRWLIk5kbsbOBTkgO38TG61tWj8tAK7bWk6UNrI+/krI+Nx9c0ISP89Iyu
roctO4AmAloaN6dhMRkrdD0i9rnmlLPdXLQIEJReNgDm9GhlUxvgGG89h4OiP1wX
mBpz/YcdaAIsqHthvForkI4bZKmBlyHeNRZ0rNvB+sMs9GjdJzMcZX7c/aognXP7
CHXx0xg+4pGS0fw9x7j0NTixFQ+gLx3ulEMv/SREa+6MPvLB0KChh+anKQgIzdoT
B8+q6pZpOS/eTtvIKn17PIcVPEnNpTgP63zzyXbb8uz22yJZR9OlMJhvoSlyIjA6
h0go84AEnIxDczqDCJ2goCXYaBJyA+KC22ZTJesTYTZ/5C0DDj0bww63PJoam4TQ
76vhH6v4mCDYFnSMUVRCnqqgfhs8zSQ8vYdTLuKWMhhwTx9YYXEdwRSAqLkBIo8X
I+YcO2KP366hG7Ksuz/SyZXIYwGfvgQrdCdpgmVKQ+N3rcROCadF5wZMTiOMwhN6
qhnaXYspaqTZGmeeARVDR2hkbW01tlu+9PJK9rHKdg3BHSyH+Ahrv28DhStgo26C
MaSCTIKpVA8yQT5akQ4lsCZhHx0FJaz1NAkLlGQQ5sYrV8JRHjoEeTcrDUBPSk3I
MUtCYZoW5DLigiR/T+dQckx0nXQLahyp7bSYCT/47ssEEmjq+ETFSu+oJVjHLdR8
32gaWaaAwC4Hr+cHjyXvnfNtCyliPlbkWKcE9Nn5S/CwZG1OapHXxR6X3kDdcYSC
d5e4i/CQHCUW5Sf4WaRMWu7Z1/qSslymiKeCRvA2l8zxj2CbuTzTDx4ieEUdfTfs
aKMHnTZVn+E3YnQ26GxrrXWAH1P3VV+GOlQCpob+9U9VDeuaKBPQTq5VAN4zsTT+
b2PJyKwn/bXdRaUdZ2dtDT0+EY0EOY9TC9Tt/ncjQU4+AL05UQBVgz/VFy/u+hxW
89z8itHHwlAnm+yLBWAXH8VVEejyVVmKNXikKOYheTxyivyX01QDhA3RyP1AK1BN
RX2oBtmcPSJDEJEce3RAP49wqXuSCr8dxziMU2eq7VS3VD0HgucmvkKj5x0/teeh
lCJMhZwhc1vlGWVP6VMf+lPu1dGQkFVi5jk60AMRoUmrfNmxBWuUqYW5xEPHFqeS
w6TIoJBH2wWwZrLQ/G80v0XZAX6aQUxT2aWEACPNWcyttQelBq0F1XCI9vtsNZhP
sMvhX6BRk5uESSu37xjxllIM6YpqiCKHIRgB1PDG/fP2+hLvfxHEVyi7t158hXf4
4udLero3pFBBi80+zfOW087ofrYVYtV+f7w7KbRDszEuBTa4ZvQ7l7GGnfLQuxI8
CIuP2ZLPM990PU8mWf9+KJBjVlQuRjye9OuvXtpx/A2jyxAJfEE0JHn4fId8nkVp
ETryHl1DMXfrJtWr15WQ0JfRfHJptXHLanwy1umn3ip3Kw2lSZJ37vSSG3iPBs1g
hrAtmxEuNOPPfsbVu+EA7TcdUZnIJDJ9ICS8l7LhkDdj28utFX+j/Au4FLgCu4/p
zqsDHjWAfPOYUQf9Og9KLp61d/wkgz8KYli8b4fJmpymU6RVTo3mOs6MjWib3kzc
uPuwprjQIkvNgxmYTQnUbM1XorS6BIvQwJY3vztJqqzDRgZ7v6CfFbcI50WTpiqT
l50cNXZ5gZdw/orJ6s6XRzal7BCvu3gP77wUXOuUuR1pr1r3z9zcSBfiaEasGNYh
zIzqn88yb2Pqp0JP8CCR416CXVecSPTYceL8kpAIC1aCz2X4qk1rzuY+TSvLVRrg
4pjOD32hslLVFYX8wwY6QMTGjP+67xAW9YIpb8AqECpKleBBBAaPFGD2Ve8kPOeH
6Yc46fjG3jiirnJU+NfLEyDOW9sQAX4OL8HMXsHet6GUiX5fymUt9AVNVnCMMFzV
CFz1hG8UvIMgOFw8nynhkfIYhp6B3lku8WnXDeAJGrBQw9wuXfpZT9oYCPQafKvw
r3KMgMzNeBvnppCyRdav5RQoav2QDF9noBDBY8sTPeezQVk/23pvLcRGPlQNW1Pf
uv7XqxxoCgT+MQ3ltxb5Yt2xog+pRm4mRxwCCizIem1/NSa8WGpM9zhH9h+X3UxJ
f79uULhCduZ+vuvgZOYH+y5MY8emjI68wiwusRU1pokk0Np1oGhJSympgAdyr/2l
NCWa9/7XW/ypz/jRPzRvUCYpnoMdE2YnZCibt/1Y8nS4HbHVD1tplnmSU8Dg51S3
Dnu7ezeqJ5ayMtbsuXTfD33NDSfTA7eJcDXSfkd+GFRg74J1JQCElRr6fIm6yhQ1
9SuZX4B/Lsa2jQgGjb0dEKQK6lDKnYNtHvSEU1/yYiA+NMe2TOdlY/1hIp/Q04YV
WdXYCZlBzyYDjalwLFYxckcJNKQ9T+5TME+YkenyPGeI2LS0Zt9FWk6d4b6gGh1m
eAKImeqOy/tHYKYRhC4KKTReH8fMFopCHOJPsyF/V/UZfHM+Wu0KEhY4iYscJrri
uDMimu/gdcxHdKjbSRERrEST+ZXXyvMBFOxt1H+64raPcqTJNUsSZgGbUxLQNJBF
g3xqNODQEjusc45KaWjIHCc2Fmk5Br4v6dQeLltRvtzH1NbiJvCL7cDOouu8jL3Y
2uO4kKC2vsm/bfz5xrijeK/YsNErpd2h4Mncm/Rbylkz4zqxfO8nFnMoZXhMnBAB
YQApB9Xh4pWUzxvItictWofr58gAO6h+yp2Ww8+R1QquMkFqdha8q+C/h6kkrjSP
XI0nKViPGjBoqSVGhQ/ppOi94LjlBYHYV5ZFeMmL9x8wFxm330UroNlQ8cUBOOWM
9MiH5xoQcdkbWH3fWyE02KbcykaiadcLeewVIEwix/n0ZdsO+Owa1Hp1K3Fal5Rs
kQdxmcOUstXrLr29WE0CNLWFi8FKOCT2u6hJW9cD9QVKt23PMggPKxT1OA0i5Tyq
Tc3ooFTc0OXXj6yOF2tNKmMkM3xirNMJhyG1i89nSb/2q1mylUGz9N/ijL14bYG/
c98/URnOl9qTLK/SnQaZKas2v89OJ1tB11TKN9Q0DUDkDh5vmRqCSmXl8gcD+aEG
UXXrrHpDFHlJbeZkhsSD4gaBTea5DLK+siGf00MLZ2wcHZfyAJF09jXWCNqfAz+u
I4oUcva+4ZEwVAgEQZGQ3GMigixp7iZmKjGIRH1J3A3I3Kv+oADcxKmX2l+MyeJ9
QjVbwlg8gDrtJ64H/LW2sE4WFGr4CTw+/e8xJZ5Yt+Ok7qZuguCOBsm9zLSd0LCl
CLK9f0620YA3AL95DWlbCMy2YJB0Lm3/6/6xXZOrcmYuPDFMS6Jy4mebHQeSx70Q
lKHibTHtgbVOlXcyYxApgMCRH7GmhyYsA1gxbTNyC/QlFjyzQwL4V3Gdd5qWRdJH
MNT1pjAemHVCwyAeaiNj/NpQbQf/SunLsXWFrWj77GMt4IlfqBAHKKq1OP11o2tQ
3huXepUTkyp1HCQlnEIIHeD5ng6Wike8S/TQiZn3SGlfPsObolJ2Bxbwc88Nfc/I
PlpZFynCTJzhC7Cf+f8WH5UF4iB7P1BjGxFQmyB4uAi82pxK3pxr6knDmcw1lbTx
hl1mxvF80whAn71MxlQUGkJvT4kFqOQNq2h6B5cWKamPBFslkDsP+ADAl1/aQhY3
W3tR7/pIeVUv5doQEKWaRIdYk1YugDXyVDfUz9drEE07ibAtcQruFerYSdAq/vhY
v1gm7+GhaaquGKM51AVTbBfcIqDBXVLXRjRwinRuanH8j00uzmMXd3bFjdfB1r/q
2LIWtZdcveqXc/fI0WaOrdrCVSF6eqDKrxa2ylZP3v27lrKSAYubtex1Cg4D2XoZ
4cu+TIB3vib/8vOSRdN7pQwC2sZE5UCrtLSF+ps0jAD9//QU4N+mMlolnLqkuSzV
Wu+AIKp0bVAWkW5MratlD8l0k+0Pb5ObbmfSsunVuHBnpxk6oJHc5qQcelwDYhNY
RUBnKq1utq9zaKcCWAaheQOycpoyJf2T8/CG1ZmC8NqwqYB7lgvQByr8jIFmYRwI
nR5tjbU4YS0MApgSYdMdqi1vcKkynIntROX769737V1tRJsegkxh7LUBrWauqMjl
bVWoXbSZQfu9ww748e5/AGyBIympgLXpw96oAMJCUX1fuMcVd9HLdRMlo+uut1CU
ZyxFuSsN6VEHcigXo6s+d5em5/GGR8kQH/yynSuLblp8z8CEsz/LAOtth3EYDjw4
7fvmFPoO4EyNM08UmT+Y+IrA62MLIRrzN/PLMm/YTTuC2k1eijJDCE8h+jIUJiU+
QR0caiDm21LsGfgA0JD1Qu/n2bNxZsF9m6yt+aPoNs2FKfS2/qNloX+GJ9AoS1j6
6Hf7brUJlhP5mGGeq/nuo6i+bKCBixql4mZJFlOebDW2vbLK5/OUR0+PrbPVDNMH
oIMZqP+PLrRB8WcyNzB/AD42EUvsTk+RQEIL9N3kv+jnKU9t7LqT73HZuWWlWaQl
mRam1zyw2cVqFF9Li+4+qRAY76hylIDMRyTgXMz0RlCdIQWOmGuvNwY7KBV7vXVB
M4gts4HO1GSIdqjLRntpHeyLIaJn97RXUCCEVoQhZHNVUuCQr8nZ29MjyJPkj7UM
HsvngXkEF1mqMtNRSus5J0Ap8ifmRsNyppyFxgreVFUXGAR8ag6hBYeOanWfCvmW
TALjOGdNehy7/3P5o7AgWY3eTMLx4Z+t1+USDDFK4Xb+KSAfQBucaG7T8jIvuQdL
8vWq7DFQRJeWtQc0F+zFQZenLF/do9h8xmFUYH0PKxyICcSNXrGu3OUfeJODBn1H
1f9fyYGCgYAxTBlJ09U4OzSYDhu4UblM1Uj4Tbkk2Qce61m2WsD1Oo4KDEzv7Oyn
0+irdKyIT0DlzVGkj+kfbjhGTcWuVwdh9kVF96U3Gi0Ywx17r0Huzu2VScAvKxl0
Y4lIoMNZ85rxCTVdqc25BeZW3ZbaDti+wR6TxwUQ55+vZQE18F03IPBjKzYsvCP0
XRIeCcMpq/RK4iGNaUXDDs6vT10F896jqtKP6/RUdTo69L7wlBPwUHqXIEZJbCNC
8WMfW/xR1AYc3vCvYNQRNnMBGH99mokbvH6RWvrulCYxLe7ele2ZpSTan+y5J0ri
WzF2h/tv8SVjTEIpqgz+sFjPj932YKYPRwLPeAZbGqF04LcwS81SnEpd3lGR3yHf
fCB2l7byIRhEG6Y+F/R9irC2Fd5RKms8sE/B7HJSk7UGCawBpzA4l0GREgzatLiG
81H/CaplGQe4LYdtronlK+I0SQ7G4ZBDvaqY6QlewnqkH9D8AwCPCtvl87RRMV6C
lfxbVX8SqXKGp6mVzw2w97qDrJLj3TQv3ZPB1QifoS0v4DaQHOZ+Sz66jsQgdCWQ
7d/8iOHwRITArzroJGOFnaqVzh125Fw54Y9exONJBcCPWx6Nu3vke+l5JXbfzeJA
KfItFoHhm/n21RN9PLuKPZ5snHCtdLIOBSsVS/sBPXVmdL1ivOsi+m+LCGnR62Eg
cHEe1AU8iQsSFDjOj/wRaUEbK23elUyblHcABtKgcG4+6+TndWnV9RUcPUfMUZwD
Q8mEDT7hk7XZ962R2TdLdXpR9bKNBT0njoTfT1nyFafZGupRZRWanzDnbiS5cvqp
E246ZjE/u4hJ0iq1SFh+8KI/DqAw5eRIUpS5JkRcuKH2DGox3icACLKoYdi/mwfA
zdfqaHdaGZeA7r+bEtrSaTqcK5/Q+TY9ZR70C7dfmJWXlB29av2waO/4mPiHNBLB
CUfwQlchRao4UcfnS8o+u44J4MD+MQEJ/IV7C7r41FIT0jBIuoxgjhw65wVCd+1b
MeT6PSSTnoc6LXlcBfCngK1upvNFWuaIhasxleMH4XO1TTtA7ft2CZq/7h4zwrv1
k4bNovVvqH5JqBiZON0LM0d2GzZWOFSjIbw9xoDHh1sFq4jU5XgoaIN6+tkd9e27
x7tKe/HaXwDftLba8in3P9wok5rJLSkrtGBYzkK02fY4KU1IMiTbY4QoT1iVdVDg
tipC37UNN7MNyNIq5b9h90Hm7oQEGaH1UJ/d1DqY9j114iPB5cNUZ9PJBehfrINu
MxmwgnKH2dCPaTmpcqD8OHdgwkDDGBucPn6aKfxqOeZhGsg841aZhAXG2xjPcIg0
4gC1k25QAtKtVxaKtmHq/BTx1+8K0lbArSQx9HyBLNeSA55bqIRsJj7xjiuGPTjw
x8olr8kv94wgZFPVl004TWSOvqY8At3I6P9k2ytgAFxvc8HZDJaviUnAHcClaxpn
SNtbiHeyxxmcwt2lDgTqUk/mlrE6E5wyx7REhlUXIf8a8GpM2fdxHpxPkqPcC6cq
Mmq7CBTycGi2I8/cws1+4q5G9gyIwgxy8maiHB6ZPV2wHRYW/cmQZLgIYVbc0vYf
74dZKwd48ClughlWLIqur8jN3hQkAK/FJ+sjHslMjc7eNa4GTxeLiucAIMlIDSGL
YMNVaG6WsTP6er/jO0aWha9xe7yvL7DPUhhIZCx4Tkj8Pz6iubouc6NyzkcWD2aG
azidnK1k6cbuz23IZuejyvTmsW5rO7uaO9zkNJBpIQIuLOgaFXQnI4OwvNDgUriX
JaXw7wlRaczjJJSfXMHdddIdhqYu+vmhsFAxxzCdLFAg8O5HzkgD1r/SCwt+nxNC
HztX28wsiNojC5WjRJ04KuGiWgiFIXtGxDqs56/Anu6MF5c/7HfULRPpWIlxBD84
JiT/lIuawKk0FEJehx3Wuthyg+kmTe+iKMohw0krmDi3nvjRylPBGFSDckmbadxR
ulTPIWmhoQbcYfDV2Qr+tzhq3dNoH6A7kZpJygwM8sKg5s0qLPHMP5OLj6OIcOJY
RJcF8JU2fqMxg/mQ1eGMRYHiWQ5+6biqDtXt1mvDYxjsxlVy0xPHHc+aPV4FxzQ7
rI5vj7J6Q5f8Mw7BwSwUdhkkc755iI3kxHJ63+YFwzEA5KTlgtsvVG9qaXzIiOiN
jCxlUBOq16Nq+iTAJFf60WC8HAsg/HP1UpyftL7OieH3rSCKTNv2bzlDtzOC/Ny9
GKg0P0N50tf+aJ8LEuKf4FMDEV0DIDPOy7trT8dtC1eA6Wc78cCchnfb7W++ZsmJ
FM2fliqHpEAI8ewdZD0NwewJEr6/pl+5+nwRQ3l/zJ//o5HXbl25IsqiimoEN/BR
clf6whbTtYzFP5BT1TlhkpYjSdDI8emO7/FONt2HJnUtajjC9dhPqxpkiRufVFyw
DyNmpyBq2PFQrKPeOj7vQLtYcoRapKAZjvZ5KexJj7Q2t7XTLl5jwoVHknQAGqd4
isBoU4KUITyQrblccFUCch0W/T+lIaBgDUXBQgi0+A3DWZNUWvHXpfM8kEkN1GF0
NZBv6K1/JN5FyXj/2/dmNzx2DpEnWSmnHi+MwTllDLgi5KiLBTTveR7mDzVFcGFv
846jJbS23wyX3dAL/AqlOq2dWdzuKA2zSPk+WLRDTK3TnV6OsPUgG57N4SZlNgj6
mGUrRkdWi1Gt1WSFf5uvvtcUiVvrdVNAfL3e4D6uf4P7vSiG3wHeFXT2JPnffrKL
utoDgV4mB8v1k6z1rnY5dnMi+wHaxOz0dLIJ/mi3zxgCjQ80pj+LLDIBY+JA0jjb
qUUxFgKugg+wGiRkTY7S9Kva/2ot++H25mVdNKZMrYRbacMsnY4hhQktWSPD0uE/
bsAae8uGfzlDBtKnKBVwpRozNxAu9LJc+sLRXe7M8pEwya9gyXxxs5wdIiv5mbGr
CP5hgr20zEcJzBBcArBpz5ZTEwSJk8iUXixLZa2btmIjUDe+SXo1WWs/7IDLY2iK
msUZkWbRrPykwiGOpYg0xyaDUb/ZREf5lmCFeyU7D40bekscLtoAeYTvmMADH4uL
SHVS0bSyh+v5pin8z4X0Ax+j4qDU+5nSJEFbOs8kc6y41nQGkDeyjX/6YBrj6wl9
f78yt0FGs0mvk2CFJNckOtvA0I/efN0SDXAvIkill782E3EOvJ7Uf12cO7zk0EoN
sIwp9KRpF0m+mjVVDa7kH98Cp3Vb+p7mpQVhsANQjJoy49Qs0mzaz84KTCUehxse
FKNOY8j1GAghbfACc1360hcIvmvEgtZgOhL7o2XhQ2OEpPOfjbPXb6Cx0oGZleDi
6ofEnuj8ePRRJ5iQmjzncwBycNppxG/kiZ5D4BNn4ihyEgljoWIuUjaOtkkt78CD
Lft0JkHwQKO7KRgQAok8Hfp8zLeZ7iN30sVsgORz5XLYrcl+3Izp0Nlh6ZNg1nGr
6eQyzTebAdnWdoY60sDDj2WNR0IYRCG701d7aiU8JPQ9kQuDEcpaT80Hx0HQyStb
5qKmYDMDHl6fipJI9ObIO+cS8A5nF5QYhE+sT++PnDlQkPpDDe0FnqF6tnluCVO1
DAy7QDkNmOeaqCuo4xXSbcqLAAsTmaPZZi4b893ugS8Rqn6iOV/ecbJmjyGz+I8o
hFrQvfeSdPMGzvkH+S7IqU42hOS7OmS/pgKcnx9JCEJ1Akpj+Tzbl+juahskj7nt
jI22bq/hhEgXdZRQIbjR0b5/KkA0glm2avELkpXRk8WB17oS9v3/9W9ysYHCQ3C7
PBYeL2vgqsQEBabco+pd29/4nOwUPH0L0vRdOTEZpzZf32F4caMMRkcghACCDOIn
iofui3YomXcDcqXNoEiL+kgzvHYKV5UGQPAw7tGrRy85uJnGtoo2BnukezQ/iyTF
QJIhI5k+gIZaf4ALtOgqxSI1WHyG6IuIeGbmvmk0OArJ+2+oaieH+tqsZoSpN7uX
0ftQIo6c37+bzwd2Q++8juFXI6VyjgdlUH7yOSJvGJptGIF2lIQNpXQWVGrebQ7f
3ragz+aaJCkEC8AjUjxry6+Luu4tQnXcOKT+4o6St870EZ9dOLroJ5IZ0KZ3NB0W
PIZCU1wFPZDdgYdXVZkU16hINpMK1jF2rprVHvbOfCj0K/sBDdUH9jTy+X42TPas
hNgwcXM8oWR+/l1Ata51muCvf1utyP+5IDdw8p+YNJFzYhLUz9OAFQ1gwX4c3J/w
ILcn4dhc6Ot9sbkd6l5rBS3UG4WqwICvyi9ken8n6n0INq3xkMJqUNbtvaE40IYf
ufzVln8UASF5UvFbsJEybYYGfAD/eisbPHd/6A+9riT8wUkWo3NzIBx9AEYEek5A
WcyzdV/LAR9BnRvrKbjekqoNPieOGV6u26XUZSp+UUEjwiI/BAFlcYpEb8JMclfW
LowLneHsofAY1mcKKECJqzZiMDdm3XIETaxDq46EogrbJAXgXi+HVZvjjlTtLGca
Nn1E0nomaOf7SavolA+FDoWfzASAKitmWEguKZNz4cIdZfIztIh6hPAmynjeNl1O
/y+6BEmtRuTfopN0oGVGlAgYEZ1PqnQtUA5SX8F2jZiAWBvEbOlGbo57wjsljU2v
9AqhpZikQhisFeYUU9l0+P7x8S6Iios8aiRhiJLNQ38LuvXPZmK4PmpgfSFpj0Zc
iXbGpzmjkeGhvxFnjoGnO/6PIQU34atFz71FU6v+7GwltItK3R03gOFmTFQT2Jz/
vtj3KdTrRv8b8NxnvIHcGn0/0iz7kYkouCO5tuYp/EGW3dC7eQvtjK+FkJTXJQo1
LDUaiMahbL4uRFzFXv8ojyqgCeqAxPLWJNjDMVH3bC49r0hVim/18lp1xWzuKkVB
xY0cSGYicYmZrsRsa+tToM0bgq5fJNxLORwcrIyz96DKfxPizC6eNxWiJxVtPFOq
q+wAR2A39mTDPZueLJRNLc0EodHsUlvBPWbUAdHrL9LhPInTzyapUlgb93wt+5mk
j3OU4V762lrM3xzLvut7iTIferWwqCqQhoGwElUHsxPGk9qZnrM1G/w5zs3yTfXy
CjaHn7REa1bLE2EvJ/6C5R8AQtlFLV8RjCz3iPOtq5WYiAQwaD06p4aIi62KGBjj
ofl89cMZ6cLR1p4TbSWQVGqVbTmjpes8raDd1xdAQ6cNcTuMf/f4KhMPmak1l02S
w6pGOXH7wCNW1pXBpRibsMOYN7LQg3Z5ki/TrI840H5cgeBFmlDoaoxIgOv+NF1U
OKKpFJQdeD8W8qla+YXlygrrPcOcHqPJnVpQh8ByYNRfAm9+qfieWyY60uvOg7LI
IPqn9JVuy63R0SvWtmtfZNxF4uz/h9aKEoV3+myj9ukqpjccJavBl958TceRsbMm
XIymPCwIPk3W5sQ42EL0T8Lhaz3onzHQ2MvT4guR/JEBRLka2gGRaXuR2l3P2FSE
CKxiBWl/0VTlHsgIBcvsTgaB+Dp225qXCWo7sOei7Wku9Z/iABOG5MFCGQSA8bXk
SFKQkRT6WHwcz/jcIXmbLD3zCBigXlsxqCupuK5LtuQJA1SWNvX5STOeB51kX8Tb
F9/j7hCVEkDwqaWz7NK7RjXz3YuLwoZ0MORCc8asUxxfaqfh3Qg3maw452lquIei
l2N/LjGZNvxDh74FGzq/j/BlIhWKs2lxjWSA0wV7s/wJz7OfQcDOAv4d+RvChQDs
ZQ+TdOVe9+ZGSIsRVQTVqS6+a1JFKzMBrd5XNJ71qxcpGgUNsOZpaOC85YKFJXDi
p4qtomB0w6Qcld1XrEa+sr6gefhUj0eBYGEtvflanyoB1a8XEeOh+UMuamuFvBKg
v4sHR1zss+TnMPrjg16cZHogrPpT2tiHM/FePZ/LZvoxaU93sTHIgpRfRPNIYGIs
Td78Xn+ZkjjhucmODIwA3HNoyj374yKgVTqe8BtNPkQRpVvJPmlkrfwxHP+VRtTq
06G6HlymuxPp7vUfgQtSgrPlpnJK0m3zdLQ1w1ai3EZcLZLt2xU0CmYh7h4i4Vq2
ZYf/F4KbwtJZdK2m0HNdIQe5huHjchqzrB2Rq3QvptutrLxOmn0+OAjwrwjLR/bJ
Mm1uKIeeIXYl4ITMx7Ek6VZMQCbV2rp12nFtYw7a80pVDejj52NweoNaZTi2nRBl
L7nf14nA248g+Nf8RrJykOc3ASBFPgbXvKMgS3vDaqWN9pwsZktfpXZRqF5yMPLW
/mxF4CXkVqTcvaS1aFHsFsg5Dgeu1kT8SSvz1qK1pH8tpT1Mc2l1I/+tghfGESzo
dO46OMZMaGEkydek/dLWwLhbC85HsSuGfZoXnyzKQG1+s9XsUtB8jHWKx7YElxZN
JlwZopNfs/mfVjlcmrMrnHT6Vak6fuchA/8/VekS7JvA0fEhPetBeSQsB2uWrEr5
M49AfEKn6UbjDrCeHyDTUYZwFkPf2hSI6luCiYBR30QttG/Mri7mVUcMAIPcolY7
NI6Bg6uzCVSx3mEnEDvrBdBHDjODIw752Sg8n7QAnYqsTIA7g/FQTtoHtN9d7/OO
Zvq937fDtgMzMesKSDPMBUg0SDYac2nt103P+k+lzPM0e5VW4XlrOpdyktRXRSOA
8n+/Td27ESXkJAN5TRNvi9A+F9Dq8EdGHRktf68tddvssmqOiLsYtPhfBOYR0fFF
4JZQ7eOPp0MFqMNIAsE8mpnLNzGjD8h/ReFDIr0cqmPWo15RJwQP6pm0B3a1AGWY
a5Ufib364by4qH+8r+fNYzqDjOjKo9srJzlHvZrNWwsCb8/aSb5JHaM4TXg7iSrn
bKNsbfBwYTL77bbaXAaRuTgdSwCI+2wlxJUBtGWEL3hKnkN+h30nM04gbeYu4Bi3
GByzsCUB0aHTssEfy1NoZ+o+38thT8dhOaKLDBFWLV65jZb/+W/Yfb+/ab/79R94
kA0I90emHvDSgrs5To/sLpKXpXrHdnGVAzTCgr7A37oLq+mkPFEfa6PhpILosXou
be4H0pcr/7Ynpx2FxSChTzmNMe56PH9DwcyxiB9y2YRYbIOX3KrXq8P4vfThYIMy
YO5lRYediDp0sf1/Jx4rKbueYo2+Xxpq3U+eUDBV8jYmdBtVKc7R6n+r4MitWX6U
NiM4tuyGSLW7uiy6g/4AXZbzn0nOnC+ci5T0ttBhScVcmNQPDYZcGqs/gfS3Wg7f
KUIuzKN8gVaEKctFtMJftjMkJZE+FD2SdiDI/0fojwiojT0Bik8Yul8aBa/ePjrT
53SEVMseY6uxb+5qgl19Ks8hEC6BmOBJUexHQS/ohBy6X++OVaiCTsqzzVQYkVy8
O7P3ZILTSGdO8Li0goJk8E5mcaZsZ5WWGgYZaqfrk80sAeeo8HX1xugdgCiaf1ez
Egipr4AIuX3YqUo+7UxxynfVIcTMo7CU5rIF2NvTvR4amm0zg4YPv1LYjkyWIdBR
pAHjNcakf8rpIMklIWSKXL7aalRuBX+JxwWGf5FAj1tDd0DjpKhPn1ABiya3VA0S
BSkvdP/mRiSjHJ7oyUxECeOZ5L/+hOAo8D+aFZgWm7ei/RoYh+DkTH9mqu1nA+mD
1jZJnWKPXFRPwUMNlMpigecRRa+Zl8ni3KtcD+9DEtJlBoD/I4pDQEc/MWCO6opB
3mhHho/T1MppqbmKGztdXd95VAohCueOV9p1IkXrKsE1AkpIVSZjNyCIUuX0dnen
GLPN8h6BDLb/b99pUn1u+iUv0/ECniVpSHNn2zUQSfdGATrNOdDLJHoPfRYyWJgm
ibnyEiKdI6mey+UDHUXZoEuTV0rKDpVyN53v5CRH0Smr7lcng4mvsICJZP2cLPlA
bN5eRJJicBeLN6TEdE5COEjhigSbQcKmbfmlSU5Ks8X5FnIq0x/jSTo235/OONfT
l4btItMoQodLw66BDrLS1pK7i8Ni1vAW1X7htvDW80U0OuQTVWO3bNO/SGFfOjma
dOFBRnQ/MTbleqZbNer4eeJWclC4CjnGDfubqefGnuHFHv3bEUohc/akdl2Y4ua9
yd70hEoNMe9nQMpEWcu4uLZ8ryzDWxaLcvBwmH0dC1y32rU1M9iONGgP3kETL6hy
ewelQVTbGEFfEXyquFqRT+DrteHxs8LE2x7KDwfjUErLBllybyStHYeHFFWLEoKK
2EhIQFKAy3n0E4aXn1KCslHZyep7VybxCd6bhovXK6AQ6Btw5zSG+HDHTY9+qMjf
0sTRPbq6gft1ydLWjg3uTT4X6QqQuN9A+k262AYC05tR6d0z69/slut7BW+FV0qm
uyAJMYscet3qGjR3g9RJa73weWCuFGuRxTLkHVD6rr0p98bSiM+fPcak9Og5pemu
3GkIHXFmJISvy9HFMSqrKxqqyLNw3JfN1rzVKMzQdEH2nVupXkQsIf+MB3kZEwJP
xf+KqI8Aroi1Q5sTlWOLYTpErqC4QXFQD4kndK9AiHskZQvH3EjMOjf8lvIWTzeo
8obDIGeF0aigr+XMOgiSYMx17khQbfYqJM8tIvD4uXXzeHLslATwyuQC+3W7vfB4
x5kv710C+FjjHwFpb3HMOIszXOjEXiBWrIxDRjaRJxQkHQtwVKd4AOTuCPUvI26y
ygsPzTSHF0NCT+i/BCZaGqBd11TPlM0oVU6vl8qZ9dQWa5lfnczQUKuznmUeyebq
P0Ox+oa6jxfvRxJQTZFOpoLWAyJT0zttOJ7l5054xc3gEHPMfWh7W1pNY9QoKMfY
t1z3M2+4K+tM8E5pWhjOnU/5Xdwg1jlI0upKa96UtZbr4HZlC5kuaB4MivPPEe8D
lRuyAQls5GlZW2JRTs1es3E5fM8BR/Q78hEGfnKdmFBRHL8ySg8FpqXKe6OA50t1
GgScJBeUHhzNoJdvSJR40ABWp2+JZOjpAq/aOTn1ZPOqaMtw2K/mGkUAzzXT9+ql
T1mw51q13AFSx80ogFG1+8Kevy+07awToZbwkn3dtfj5sf9pncfRXJF3eDqqBkz9
SqHhH3LXbGS1Fz4D3YAFnIBjIjWFTlk4/kgSt4LAhB4oOcABq4pA2zp+4LQT62C/
J1RgCiTmRRuYwizS7Z8FzcQKJIsWKUqJb70P2VHJZ1WHwKsllw9xdq9im76Tq3IU
opz2uwMV078v+yj3eEcCLj/NP070ey/1G8Q22Xv3ANANwYYhXiOZY7G+5coHJX5z
DZVixQbUN1/Y+6rw3/iAoWUvEchbeq3oGUVfW5Bsidgda7O5e0XqmbhPIvznW7jd
BFEbw6pqp6MYKitZUmk5MUlY/Luk6vlqSWwn3ekkMdulOmIJ6D+nfpnbgS4+rGnE
5iOGKYTt8onDyMYJDs15WyFqTaVGsrrE1qi8wdvYLL9RNoQMLCfggEVRl7H6hUzI
gJzRMcfWdHt00jPaVic40nB96mI9YLa69YyMDhTjOhrc2pTMKk2Ame2SGQEEWRo0
Peto1AN/v8HEp8nJ39ZeVkdkfW2wetLuNZEhmrQxdt84RVOP0rtJdt8lYtG05dkb
LZCgaIAd7UJuyIsodAvo3pz6k+nwVEBbviOEOF1Vs2S4AQiai6vbQY3N/IW/muAQ
RDBuKS+sYVIFGSl87F/RogqDqX6JUA/rs1M1gUQHtPb9Qb8jXtqNeB+cE/Eonm1/
ukVhAIuQ9b09qHNOkpwIbbRdmp75SDhu3UXRILKxlCQYrtffDBjnQVg2nVTFT7fK
oGNcvFqMOrGbO+fy2lOMIqhYcmv8hhrC1CrJmmzb7wt6R2voe3eu1gGupUMeusrf
dbBNel0xZAidZ7IPw205LI3X2XBz5fGOFfvEx5UD+u1uUGN4RcDpNGqxMSFi52KC
PSkyKSV+qNdv0XuHTk7VlWcZWAdZInCwLCCKBIiGqpcFAMZZ0da/qw/+O+dWwdCE
eC5yqVAywNzPYFLBr4lcbr7ptSunEXHg642fMNbW8IWovBB3MqEaIMYluvd/m8Wy
+XWJ00ZEPEkxcSjZ2rhj+5V5M7XPfx0NLbewPwQNjS1h+iAS3y4hdsy3B9CTxFGo
HwcEtupTLdOjpQO8cP19fuXmqSirlDRAd2RSti3/9NDPu5uc04on7DAFjzURK7if
DWTzOcLz75o6PaPIvdouEcsajp+ipAuwcw1OjdUzFTF5CsmACXKctFXzSBLlgWWM
BQUO9Sftuuc5bTX7xGRkmQRVSVWZDFl7xUEcfPrrMkwkTmH8MV4+887XSRgLH2oX
g68Wgzx4x/m9TMp3l649RpdiWbdFtUMOqV2r8RIifgLc+TS/rfWRnqQdi9QLpHM+
+1/LQj1nhsvsDN/LiggoH4Gi4eTxjSIwEllE/Mm0CWDt7FtDNh5XniYe8B2HUpKT
CSUShn1vNoYtsBaxv2YOCKbtceIZWBhb+/5pkQF1Nz2/AmSlXs9VhqRKBI+GY77X
o6sFjDjHSs8Ou/PvhNjD0ekSWmFdRf530QeVzzLbGV7coV0fOkNHiDpSwqO8MMMf
TiiRSjAyFyR4otFysN+Y94gkPjAu8rMtEb11pq8AjEfPbIk+yCESb6L2KODZw/ed
UlMVwCZsjArmSMdu/D0i6WOa1iXRplS2++0SrFzl24m/VlR/thWeQT1dgl0n9H3B
bDREegHx6en0udGwBP69QE6iMcHH5PHVJeCRTA0y2PND14pmUryirXqyZiMgCaGR
j/0f07vNz5HDlJ27sBj3E5FQUQEuHGNzfVRNqITjinz2WNiDr8kfuEJyNIsYmriw
uIsg0lPqPoO0Ent408zuCGsx0IfcjNd99oKvQUm9lwSdrwwgqF4fbpR1gZemYrDj
MoLbBMVoz4P0vA25zgYa9z3vhbiPQRV1M7NIW/hMi6ZA3zJepPe6an4UpPnJNm24
cF0JlxvpHTN5TcwnxxpvdKg/vmq2d0fPBBLr0sNnMjYc9pB3VZT5agZvHvnHoEnY
cO9f0JeEXVSZwuci/9pUpBnG3HM2FyL1vd6n0wRzv27RgEdY3MZUP/oZ3QfEH5AX
ZhjqDBVquV/GPQA7LaCVLCMp8mkPVWLjq1vn+OMxEeOU5M2LCAsNmX4LxkwxU9dX
lzWuBqf44ljngBasNWiF/xr18Mqce/Hs7SZ39v45D07SihRfcA2oQzz3SbFXkDUd
HlEdcnzK+B1kC3utFTJRxycV8+9o/DT+SXJNdg8g3iEbGB1/JjHQ5ShDrLaIO5OR
+o44mROsOjYeceCxXEY5N7E5RE+qIbPW8/Vv9ybHobt9t6Xz8esiv5kTZrbKPopW
O+xH0O6nNi9GHZnGw+DuTwRcmFJVD8VDaNtR61+RaHKBkR86nwHocVgDxylj21j2
T8tGjZSlXmhJdTQ7BaOUfJI4jMq2t62NILfvc+XYJ5i6olutOSbMb+QLIzpadlZe
wo6RCHsE07qehUDF+lxK8lVPNYP45g//WYDI/3MLFF7+U8npcqEhArm651YniDb0
pGms+ONhIoVRPGcV8Y1VZOAKQ5AF4AJxjAdglBNQ5xVM2KAUPpYkycshwSZ0/8Em
oEMMqm/e9DS7KNafdIgGqkuJygz6pH69YKTXviFzhBeYYMLbwlZdsNZErd8/rUXP
6jqkqRRIQaelr4gY4fMIbqNoSVhWaErSH4LkS+iOFaXpgvxVILnS9yu/lAwmMn1K
wNMYLXTHkMpnGCcjrg7Aj63QHYCOqXL+LQ66Wv7SJZMdlsHvX1eeLavxB34iToZ2
d3EJzHym1NKNUVHTCqT3j0+YpFPwMnoVlh+oGARuqt6MgNrzGwOqcC/NehcsCI8t
Kft9GP7pZ+IaHZg4NONq6WqFrJy4j2RjQ1wQGsVqn2GUUNbhda7CHEwCq3Lm36iR
/T3x9CrhfabBgdTllXGJadj8x3pjcZuxHW1adhvG+WI5Nid29kCosBI3pRMEetAJ
9HeLUQubdGwDCeGS9YAYR1mDGwmqpYiNOfc2SS6MjXcUBPVfxIQKUJpstKSt/GaF
dq6rDaqBP514bDVWj57nZv9KFYHbusCgOz2RgMR8vG4dAim0dtSOEf0cpog81igr
662TvZKJWVIXLVTWpBf37hTR+LJuClSxq0nV//BdbbDluUau4adOiMor02T+yq4R
uwNTaqJPD3Mx4NWcerwD1EVskgx3P/X8520jqiXuiIA+r8w1oYVOgux85Yl+HMK1
rXRR/ifdFj/EU9XmRFcXza6p9qGfgH3cHvPs97K3oK4pRSrFR5pZWYCepYOKfkjM
YkrMEX9hmqU2dUOcWiGBwQUuE6y632eFDPFrpt+PoPzkd8DW3G8naYu9yEaK0KL+
Z+eW8Ks5KxFKVrVi14vgBQ+34j9+KDgNgbCf8H1OjWXY3VnSR7OUo/0B5IaSAil2
IvdY4rhbcv06I8Ngt5hnIMUZokh4kYsWsH97qgsX2ux1n8OFkVU/V8GcN8NQMxxj
JClRuL2+6dZkDbvwRJBsIPR2ZjjneBQiVTLNCDn1sYBGo5a3mAP5jCp7xljkhblV
Y+yGSpvTcVuqYm6b3ZKgPJEf5hGwQRXr1+U/v+4yNKkiDBN2tS0wwg2Cgn9LAVxW
0UdBjEYiYAvK5EQRD3xgnqRMXc3NN3E2D5P49d2vXrsBaiIKvaDm16TYHWZAom3w
A71n/eHe41GzONEuaNZ60jP03oRSJxV1kFoZfDvGrDoSHm91k2Kjc3KPwShm7UF3
kSPNXrxOJSrHW3sN74M7O/6gqHzqxiAzxU6QXDIZZMUscA3TlzN0+ushNEceNZCB
jMadwh1QnSDBJa58EVkS97+HGjBpYsV7Rs5EOECs0hCHiEp7B/36ycVtLtZ+YxY7
MboJqT1UffZ60B5DEnLKWDqGIwQdzJlbBLgXe6uOTkNe/wS2z84Gmv+Kf6kYmC69
aiUnedH4qtk/6p3aLIO5EDv8Sruug9xejCfpCwK/AtdTpn0pNB+kV7syQqiJO0D7
HE1I+yehlTHVxWZAZr4CQNHdnvl88YeaDgPhxkai5+94qaUYtmbQrzm8gWqExhUp
NSzhEPw5gMTXmkPLvPMBuOkqRRKchyiEI6WCQLLR4KqwR3PLOblFMy2va6l5w+jJ
axLctlSd9N0sr6L8tmrxFa/b1E4+viNPQER4qqnkeAdLMTs1JQ9PIyRb3pWtko9j
a6Asq8fMVFMjAnNsu/92vjU233AaFGpsg0CIKlTVe609PBpbGIQr+0GLPFFM3X2F
UxYPrGfHY9bGEMauhdaXC8bCoJtdEZE8qvCHADDnpjEl5aAlBWhXg8CFNwidwRzN
hP7nUmNEPUdOY2Y1yigDsgjbgH5gd0YsO5cvA95P7+4GapXX84/RlyXoam8GeeFN
gMaWkNAiCHHrUOIzUpgoJ/PVF11ipwCZZcTXnHhk/88s18bsEyjJt4q8hGZn4A+m
fMje3KdTQsUX6GTNwiheZkrZDu6VeuRbxb60WD5ZOJ7+iETZ3AQpg6WfIwUkAnzc
4IGcYN6fiPrd84jLoE0tBreeyRVttsfO7zEhhY8Jc93U8TW5WjsyapsLK+/RsXZ+
kqlZBVW7kCL+sJepD+ilyFNndBG7USnpbfZKYeTsUa6uYrL8P20M6JEDnxTyZn8z
dqhiExQIQPEtODxBbyepbmv9kQxPUn5+U8EqL/+hfSE8D3TjtmER8/xi82m9ou+h
czRNxhnNfLGzpudUgi/TkzPRaZAFb5Q47s0uyTpjuMl9kvxtpJrz+thTeBHFj5Oc
++vYz7kxM4N9JDYs0qt/CdXOPqZwI5EAHF3fCg08Oiwz1qmpPaEwvcdrLYfVz79l
WGVbOZvvcos6tQsERzA8H5S7aGwAxow2/VBenKfHBRdae/gaiz3oimPxTPAD/qiF
XT2sRoaNkawWKOwWBuiLMT8bBqV8y39H6s3wsn7iuS3Sw4UkiYQH36EYvJDRJfEU
PosutXA+TO3kCewRfqA2TFiNjTQ8tci7+hw2Vxu99vXdzoBzQdB7dm94+V9TyAcT
eBFrHLd6XfXjmIkgiN8o1sv2m+s4r7RhqeRwm8nFGVBgCvoWO4lQYxZtJzHLr/DW
jOqJAox0SGYWWSQihwp78rPcmb6FQnlOAvoXMi6hy92hkEDpJtWKsb7n9O+k0UcG
+rA3tG5/7C0Ngd6nWkdtIjeilYXIFKS5fjJ7dH1yklCQQHLmnSimZEQ458TOaQN/
47CI7f94hXngOiCAQDY8RCSRCVZ9dZ/6qkprjWZkucKg/ASN22VqxoHshCnM6zde
ioiFgz9dTQ5/mnaTveRusA0+ADDuPTtaIvp35Abkb4jfUohdvfLRE75gXKMMYWph
x+mpcG2guY3l3CPc69etIsdL035FdfSZi4e1s60Mv18Jg3+n3D4D4gMKFL+89ylK
rmX2YLnI11RjPjUSZgGJj9WmFiWPvtJ0HPFPlZR6zrFHxB8d/sauWBly7CovIozB
rLq3UwQMA51p+v+kpKCKpP5iJ8142oe5TfxdCda+TpyaTAE1MxxL/Dm+mF5IVWPs
eUaDCMQaVm5uj74qmOX9Nhn3IGn69neDNVg7C8ociHC7XKoUKiKsiPsmzM7xQHc9
qKcsZwRc+tPDmVe30tVwXHgIBGKYVgBBR6tEl9J9jvlNVwAf4zwvk5WIuF0AYOSQ
Us/z8tSFHHc37+b29f/0Rh9dvVuhyKnvT5T5waLX2kdSNHnzrlcbDfYuXnc6dhS/
vu1rPNfnI688OwCTjUCnH/5imOVHzud+zPfgM6z+wuXPmpLBny01hSq+A2jpJm18
g9SghKkyOTF2uuvCl169+jjYOP6Iyesv3ytOJw2RJctj60wY7YEZAS9Y7C2pxMyn
SQC54kaCxoyENDS/YEMW14qg/BIr6uWov4YggnUb9c4RLdJxgys7YZd70ybg1HHs
qDSIOqnH0LJu42pobO1weoIOb3aFZFXFi//g0FUDekWz7PzSral37W0bBVbB92dJ
cAOR0rJRtNPXo3+s4Tp4zpqC0NdxiE4jWIX367B9LqPuJAQqhcJObLlppIbPtabT
P6QM7075YwLT3Fo4O0w9z2CLivMN+wxrklHVNf93dOo7RR8XHkbD9cB3CfTex9Fi
7tjVm6Y3piXMRyyr+kIOujdBgxrlrgyD3M77ntCZcAEEfDLYG/P9mxzlZu+5N7xn
yFtFi1j20dqH9Et2nJd4ukWIsWtFoH/SSQOeT5N323fqV0/XZvp1/SL8+CNEKA1W
DgPmObbOZX4JbaWUCr9ppDu/a+BwdlKBJlC3gkcrF6lEvYD0hRyI+9hT73XqMGnJ
ryipuFO/kbM9WGsbT1t06g1rDSq/y4tEgM09atFWlyehxL8C4BM4rSnlr21jyHFq
jUd0pU6HhhvkvAQwozxr3zqIZKvgbI0GbLS6IsOKaZDbYumGpCROnW8L17ujby/M
/qeYvDK9ofQEFeRrQ3BOLEdm2k1G7yp1Bxct0dZ2X9dfy/M7Mnm6woT2X/v3+TdE
02/2+/s86qiuVd//2OSifvj7H35Zunk5a9dIAvBRCEdYQ+NI0kiavncMH3HzQ8/x
RsyFOCVe+OJKmD2N27jrnqSZxrs1K3iLwQhk//rz9yHBLFZtJzQJE8uIXxMBt4ph
1JYx0GXWtbqY0C2x4yz5T8CwnWLCSt8pBR+aPMMrglT1feUPE8FfNbQYacET/XH1
WBgZxfh3Fmc8HbL6M+TjNCKLzR3ZyCJe8pRRBVI7sHwsJAhjp54bEZmyqeGZbpPu
UG4dYVPIZXpRHMOAilMab7iX1zI4eu8KAa3F3wQDELYceMs3bOfww+6US9/PZQEb
mizBNGPLspe0Ie71eqXW24IC1EajSWimdWdKhr4UL/3o6uv3As+xMSNxgEGfUOQC
nmXsqtapKWhn1YDfgwjfSTt2x2OJrnV9ByPvzdWvTwOlICIwI9wRZDLZGB7HcvdG
QduYCCOHV654Uw8Wqifg/thEnO1EeJSudwdLj8XO9OM3Jey/2iIljgrRjkeKx7Kg
2f72rgoX3nYWwDD3shQrwImE5jvaUV9KSf2VZu99u8Q2ZK8f83U4gKW3la5dxUS2
LrbkqvgmKR2j5raC3/SMJvOKjPTNWh6qibwhzKy0RZzbLbuVnjtJ9HOdTfYc1cve
ozJUp6LSuujRV909nWh+dM+b55xBel/GESJ0XVHkf5Xod9dVUgyk7NaTOYlKNB2L
8+7wG5ZRSSFFsek9tumuSoDxu4eOCrwsb04FPR9RAGssL9iG4dVJJlsFygkHstnE
9ebC6zQFPdCmXNGDQbd3R+I8APvUHKItrIjPdQOawIUwu7JurKYOB6JHCVK2oQQJ
/GIRbfa2AGV1NZ7AydeVdviL9L2HTwSr1X4eD3RfR+tH1NkpNe5TRocwIYvTeOxd
YgCFoALufFvDX83nx1Z6TR0HCmZsUMCKAiEkOYurkoiPHmGVfC8VBSHr4kYvsQyr
QFQxPH43frp40gQHzfJ2902k1GF45wDZhgAI7iKZILzGiiww2zDd1+1dn4d2INEh
ErOUMSPNX2GaI1vqa4lGMREZzbHGObiFiau09ObvgggaH2RbLnWPy/EitAH2p0wf
qOx0TxeYll8HxCBSJ9tKV9659fBf8ua2X+8v49nA6mGYQHDWZcdZlm9OL0/HmaUg
ldvIE8asiaTjkhTKn2G9R8ZPae1snvXs1X/SAx47Od2kMzDmRqB0ynJv89gEB804
btBtdsPXwi4x/uaps0U8WecGzgBq32quTgDWMe5VpSOkWB50RyjN45u2L/YGMy1f
8Gvsbcct1iiUm6Soia54EnqfVQOMWk/Vm9mS61R+Ai/JzwDHqO7uxqvdFyOPVw2m
msHUEzRONdkptWyriRD9k1fOQ6V5WIybVoGa21qlvPapP197qM2RRgcZyt3W/tPq
uy2cSPnf7aJWUagP6YU1zJspQqriNAkASJrF8Iu9tl/21Ccg1HCwXPO9uoT8Yu/r
kMVTRKP8/DPqpidT38HwL4jircDv6vPRuWtt0DQiWsMhkRdXumOrVCiHMcJbXoZE
D5hNslG+f0oyz0tQwIRT4Js9r2JAJgDSu0A7s5KNKzXpERlOLmk7JuTb/b1oibuw
JS/7HJe70NxsoCmpIZ6Ecy3kxHc6mZKstL5uVdLgF7sBJsxnzJra0BJqkRAhXqX+
ntxsM7OwhSFz+PlXT35/GQPfItqvz8eYx0tgYeqQ0Gff4LM7w34ZY6tlIAwqITMG
2PtE9+3PqfaHBO1nuwjPz5NPHYQUqS7hHthiuMgXyM2wAT+p97EMkfnvqnysLST6
Kj+G8//t2x5xiw1tWDmnk3yWqdqham6r2fVm/lWuRFIWC+63NF2xobuIAZo3dIdo
EzlGE0VAfWYd0OiGYfJ+3LoJlAUHzqS8APnKaWE9PTqYtmhlePJQ9H/uBIrVZJ6g
cbJc8joeQRZqoIHyddtNoLjrVN3bbJI9SGK2isUSNkHRQPdcOoc0T4Vjx6erSuQF
R3Ci9/GSTIBmL9pW9dFF4PwaZmwtjDkJuW0YvsQWHQ4FBeMBZQp1xNNramBgVogp
aLxScuse8SO+bZDAjJOAxzWHmh3p2CeSiqH66B6q/WvJvg0U8pXNMZu3lIvKdHZw
Ol8fQfi/g7bsZBaZ0wlc/rCYs3NsYXXoIhAnu6GREsPAYNfRol0JSdd8VDlOFoPm
sMq5FVIvsTYOENWto+K8R2nYvKJoKY0OG4tEj+FC0ajxj2tw3CveTy8SnuF2oKf2
/NdI9UDypwWydG7exTWJRtZ3qdR5KvwllB95rEqbekYXSnf9u4h6kcUT+V+L11Ru
h4o1LZiFXaeoTx9i1kirI3UeG3K+kka+AJJ2gF08kTR2nKCzMvgcNFG5PAZ4EDsl
+Rt4vj0kq3AvEXjr9ylCkSDdOZKTTuBHE+4W6nMlH+xxbGYrAnNFuX2n0AQC4GnW
339GMn+AXBPnaBdJPppufsYgG859W8/fYnqkG/lxwaD1wa7RLJE1dUChOntMIITm
c1HyR7+19wFA6UDRTRGVJt40Cptz3tnmNzRjYUAuvJRKj4dJe/L9yDFjhwZCGTzJ
RRevk8FoKTVI98OoVPXHl84D/veG2i9z3cy6rE/lVdVL3ph+6CdyUgQChzXc6JEr
CyojuDSCpkoeyzfrojJqY8MZlyDcc2pww8XD074pK7lt4Ij10wVd+1UkZSb8lEUx
8viXhCorkx8aq/jkD6kNAdmnYWvU5EtwlIynoZUkaEAxa6EifuObdRG7OS3sJRka
1m7qkRKkhzHu5taSmBb3n+3aGskPXnwHdBz0W9XHMbTbxn92ojffPiQkqE1d4ZgQ
vrfrgGct3WG5/34wZVrS3xz69YrsqqMNcN93WK9MVijvm0H9r2MnIZP93X07rQHp
V5hdca4QP8JujlYAanBlNQqOPjsn4nOUnzp7mP8WHRyZSLdkhpn0OzNRmqRh8G1F
GOq00EM62bsidq24ezXUhVCdYE9CaSa+INSQvQNAmU5YjehZ3ODafF8DQtHq5bAk
b7Via12Bn78O8VhfhhH2kiKfyRHKt2o55kDIH1m+PLfaTI/rQNMMbYyM7UEjKF/b
bBA6aLNNyg8u+FDxpR7oLCGrsDVKxELr7MxEoh9EzDKWSFJ/UUJH9i4ec9XQsfOj
5M23IeQSPMqdFsEYTiwhKsmc1FEsCTLijKTvKhYv00HA9cKTFHt2zOywWk212+EH
OFLqHc5zHYXMPVdQf4VcorNWRnvDC8OH1iv4WbJzOeL93mY77nsjoqs3VlOjc09J
EX9Wh0gQvzph3iD7qqyDL0GoUgyuJk1kp3FOg9uUZ5S7C+WJ9RtDmcKBdtSk553Z
kH3Z7e4A7qv/E/cN3l0lQ75nAZzSkRgD9sawx0G51meyP5BWewh7s9kUH1Ha0j9Y
hIlC7GQhtW6ukaKRnzyYn7Qr4/v9hQrtrmmudLkk0mCydyPY7OLD92q9H4I4WYzo
z30FVMvyL+sYQkpabBovNg1FrV1vDqh5hIudrmbYD/GHzJTG0+P7raTJTYb5xHuc
x49aLv2Y02v3NuRpEEEqK2coxYU8+o5NhFi15ssT+0G0hF5JOEvkTEYVDV05eRV7
i6B0KUtVPE9XkzjOi9q7HKvnrFnJcRcpPh9tYypz0uVE4j5axQQbLzYoEXwYyg9h
jPu2fwzga1zZU7DULiV365a7djz9lr+3hSEV51kPLYd2Kof6VJX5qhgg9OSACnk0
MTtaxSe+vDjkKIfvzxuNbQNWEKNKaqHMy8O1HtuyMeBywm5iKElzkwW+xhQ1fVRz
P6bSkmaIHF6ZeXLjg/ppTiToBzNAPYWVlP40C594D3GQmNGti8c696OtfxjS37Sn
rom5sNqHDYgez2rENpadr2JxzLpWF61yN0iiQWeZNOlRihvt307rPhxWRwzJBYCg
T886QAWphtlA5EQ0/zTr7w7zj840inBuY6F76Meh8BPumjlyFmFGb5s6wwLfdaLR
hg/OruESRtByqwoLClpxP6+8uKUw+DenrnhUxevcGdroC/uXjWvP+zbHXIX4nfFl
/zJ6423aUbS6+hBvJ/OIAJeEP8MB7b5yFZiFecgUZ11bN9nuYEkYQP+efhBkQSnz
XhugSFE55PT72rqUT5gTE3KfXTC5cHgnvNmrd5zsqqjBgwFvqVrB76vHqmv2YK0W
TSboigH75cwkzzoA8w5j47zCCpKH/0Dl+FvZJCJBLEA3JC5lNRbRsbX6Pr36Tbnt
sH0Z5ZEWZB8POaOw/qBHsEndXlWEow4VjWvic4b/weijzoz9IN7JmcjMxTpnCJUN
XGJ7wBC6IW4ZvTYN7eLhJvC8txdEFIVQAsHrnS8Ozeru6/FHRqI8FFIU7PPGZG9i
L7yZuwFxYVgV9fc0IlU4i4PKYmmdxu2hAbsugN4wmQzQnnGbRDNhWvGFLLNfQPfE
mli65opHVUm0i0ZHKgN0BnqiaD9MtLXtxDZtdoRLsUjQodme0UPsLJUcJ/ip0H9D
+g90i7o+B7YDqdA0y8VoaFoza2w051FuXNstk4+1IazRgAbIRgQrjE2QuhchTHQd
0RsSOy5MA/CAjCsfpS11ZyxHZWaSqEeeALI2YXzRMpXJJt736QpVHjn9cdHAIGbm
0jIEamTMCudwjS5XfSWQPVzb4LrZ6mijIEOgu83uGa1PqsIBEli488cSv+Fzemwt
HMajBI1NGvgF/e0jbtnKdjOKo0w7dVn+2bWJ0Ygk115pwWUg++X6mvbtJj38FCYo
MoTN+5BbyH77sn/IN4QBaClsiBEQteS+a/YklAl+caBXDDN/8UDUCIUiaXCYxMDA
92WT0EhfOQE+A27LHih6cGf8VJy1prj/NJ1Uz01WXkT4X7td385DUR1CwnVsnjMs
NQRmhRYxyXtDDOEhZba7zUQwa1XBK/j0bA7myh160pgtT0vpS181Jqm8RbUx3IRi
KG0gt5Qll0doBtDsbcsdDGFHMG5GH/pXOeGt+vxnZlTsmYuAdpNrf3tVynug0SEK
h0lIBvq+Tdl1r3F2WBNnEb4fKGe0FGhp7M0XqS1ZQg1QEQ5wz62npSgT1qj/uJIh
Wm7HJaqACUDlPj6nggkSGS6r9tKpC9RbRpzehOvgUUWO5F3oqg9MugwOJQfcFa4J
sYO4se9B1Ch1PV9Y/hWbb7cDr7IdGhxCkRDSQONSmjH+b99T4JoxCpoQ49vzFzzv
XXlC5Xpt38hHKzN+M41KlYvFY09ZzOOLXtEnHWM1azukXkfO+6hLqN5b+fw8Yfqp
IuwIF7eJWf5QIVBb7caUElogBykrFKo3A7RW+9Xt5avCFnnta2pKWG1vdFqe8D0/
kfEh+8uQe/eIP7VzUZK0XRlwKNyGIfobaE5Qxk52mRG1qu4kUyXmVZjplbD+6srh
J68ztN+x745JTDItI1hhpxcjBEzvuTPhsHyEkzhw0lICAMvN7rGCAAeIdic+I7Px
QLgnonU4FmoUt9QRU3GDD3ebHW/vWxge23WwIcFEMkiolpkkA7RdVfcJ0WZIYJl3
ciiw7baliW17Txl4Vs62LCYVvUjeTr6uIeSnjIoZxne6Iv+Pe27OCyieFjNyP3gF
Ypuz/zbGmfIe1q2Vv/90S90bmi16u2a0RzM5vMURLVTJ13WG1FIcLSN1oh0ver/z
U7utQrTLULDI83F82/jporB9ehKpU2D/0+kNMlrqyfv5nhMMI3yg5YwnooTNZkdk
hypV/UmXveT5zuBXJoKN4wyRXbdFP56SRneb8Tpw8nvMNtpSfWUq0f6Fa6phKZiD
wVGUYW6NGwc10MUUwikNzSxiD5/H+fkjtdKXrB9D3AilMoM6+LnlHrLKj5Jay5IC
oZJ+2obzSTUkamkUUmsW3saXuwv7ogvnmvmBzze/Y3TG2qdX7AIDJsU/UgYOLNf2
Kr28sD5Ut5UjPJAU/I9eGg1r4hqxIAAPkLey5VKmaMLM9JwgKnuAS8uu0vMh+GP/
Xxr8hp4Qs8rRbDr0L0zmRkoQiUHnh2jB7DvafsAjcLNVTLnTfk6i13hEosbaHyzu
iTVhw8FfKMIkC4kIyfp8W8XUZ2s5Euk3HeR1FUfcEMuG0cB09zAd9p8wzlmLRKId
rYCrc1wQ7cZl5niwlIPFAGrAxReDTFw+rQ0hRYKw2kA1DolsVqN4/O/OHuzmhQ83
zP4x/z2JDiZb7YlRCyB8yYv4Bu0W0OdNYLXFewFvSjMmcsXTh/DloO3ev2K244wR
oBsHWzRAK0bf+sAk15IEgKtwV/B/qOowCxcgAjvKnihUaP2JGlF7c8YZE8RTfCER
u4KRTW7aPyYCefqxxhYPUu1AcT+yLpp+a45SONIuSObFCDhyFAazBqAeiAPkl4fl
DcSwapejwzHo2OSaviyJVgD0TvlOUYXnzPWE8hraStXNX03xYWsnr24q1LkHVy/N
BFGARQBHfn0U0paCUGp78mH8x0T+DvTGshVDcnC78tT/d9OLBD0ZV3wxh0wsXnXt
iAx2cF9ld93NufvEth5ArvhuzBOkX6zZH304c8ezHr/k401D5aX/xZurYjdy8Ilu
jSvhnmzxZ42YRPCsSqY4ERElYRoeEaIkztAxbj1uGuvTs07Z93OQ4bY2lIGgcHlS
RTvEMJmSr5wbT6+Ms2xXEwApfv+mClOGtu0L+vJet6EMRmRlbDR0pNRpvHbbtNe2
oqOEKhr4ulk/KMhPiR2RY8gdUlhhQ59NphpQdpr0U4ohm/y1mOu123qGOKzjJv6q
JNK4zktKr7OdnCDV12/Ookz/E3Gw77mjs8j7CHR+fsew6er1gJFTrAQZFQR5OAIn
yYWGd+AZ6Mz/45lv7pMyS7own7rPHQzw2RtneOzAmEw/u5FVpKmcvME2+U0CJEbS
/oqDCjIhWdIT4xJAdVqqNUZKM0oodh/A1yfb4Nnv2mRVZtLrCwiIFbTaeBBjhrE+
KRTbzZ9kqDkpxQ2X/g2sBai7/wHNZu7T5eRZbkGJcEnwq4kf1kFFP7N2Ew/MIJ/o
KYmePyGb3qH+OsFU9fyfT4u7YTU1C9+NzDig5OWHVWi80MYkJzTkLJhZJpPauZGT
mQhhTNtaiEjz8LGlrmltsB21Ar6OdNgSt/RXSOY7PVS4HDcg5D81o3lllu+6pjk+
OIRttltWkJ4v8yIPBeV3/nwWlNh5mH/n6anQuD5QXNI+hLXf39pdNuCHTy5GjKz0
6sP2Q3VRzcywu84hoJRP9ybFBx/T3yitMiAtGRW6YOqK+OAxiMS/+4kFh7ohqvAA
U+rYV/MArC8DTesf20VTjXJ7VpctW6rXPJV98SXFj/hZYpejqumhYWDubsRIYZo6
70AalmZoxrqfcHKzoi4Sh9vJPXrhHkTe9k2EHufgBbjdXn68HIa1uZTFf9ktVZNs
Qx74RxiE/eGY0kZ6odFSAkh5LXl/N6ZRqA00HMJspaDTeUR8yCZRl3jGYhQG+GMz
9u6sU9mzj8w3eSpx+BxxwepdiXghHFrbX1bucZtQY09GV3U8hFEf+lMfYnAPdWze
vkqqG4Zom7QQfECgIClO1sjhbGkkYp4CGNfVJhZscQlsiYCGceo5ReCzdw3JtxHq
mnys78cPe89P8GIE3BXCscLJZ0IjU4/4c/BAJJq2l3dhBdr4q/Ouv9/Cw+LN7qLI
NbELO2Pdpvv29cnFZnyh2Tae0I1ZgNwhSiFJGodIF2wJiI+JT2lWGA62p4El4cv/
c3ootQZIrL8k62ODQpxYx3uiodSSbJqZy0TQMzArodqDcmE9/MGhREUZ1zm1MjOt
MlWx9/bsT4D5/TEBubSJXAQcr1nRdJaA9gmcKRk+SY1gN15DpQb56fcGG8qC8LxC
CmvoFYtCPKHYUvh29ZqSeLcozXxcVs9n3XBKwqIorkJtMF5f0m1Tk0DopJhxGYMj
neA2sBriP9wcZbuA7OvUh7ZMJYIkycEb459R04pW18tEBDcxzkpjtjuxUneOHTcC
BIStUWH6YDhLteMtVb8u0k9Q9w6R7lFDHlWCZsl2GQmIhWjlT22KXE1iSFKDQxwx
MmKSijEbxey1VA6YkI3hcgTu99+ERud5YHiz3ndqolmZgZI58RB5F7l1JsHp+BlX
lIIe2IVFIWvBeuMY28tV760zudOTDf+Tjeu7JBCcMaFapmyw9M6OUAdGt5xV+nni
ojrYaTtgGxIGMNwwjm/UJ0fHAsatw7gImZRnulHLSUjiUZuDL10y2EIryhRPnY3a
YfpVQwqgZxtrjaJ86AO7e/IsKKZqnHSDHUDK8TZonvSMf8iI3LBHK4rGaOn0V4qC
8DtFrTGxTkGsSwQxDZIO1sMNCXVbiA6JdPJolhJ/asr9C55bwh3xnI8+jryN4GU7
UFjsKIUcDtuOOyTQuqSmK9dETwM2vJ5H7JhiB9Q1Z86qrmrj2RE5DQuDnOyd3fIB
k/AeXJCNlO36RBk9w0dJ8QAF6jHAIr4QI6vqLGSeS9ZQyciKdJ3q7z+n6o4BcZWI
WF/zd9taT1F4gXgm0enhtAgzxm6ILSv+wx913dhiUW0f1k30CcQAt2swycikau+N
RuPpMBVSaUw9G8VhQT+9ODv4tKY38dfXXq3VVTSSYT664hqbHh68UANLDLgORh2I
pNuhxbdaxTZzScxI5Gr7DGFgaz/CiUzPiNCR3ezgfBcCq6NQaAGrVjxBK68j2fTq
AhF23wIAqV4Z2MSRvoYUTyvGiHay2WCqkzr5dmpgZ6L9hRN2blOO3dAQ6GiI8QXO
cbaphHTYvoCoC3Q1Z9BcwTaLNVUeR0NE0u9eJzc2OpBiC5z5rQTTuSYb7w/UHbVA
TJfe69V8S23AIH8WRzwqsZ1xMsw2Zru08kndDuRtMmtb1vFTyCjw5aDa14TCp2ML
y+3vBMffqsKnh1wlzrENYsaz2r0aHP49Yfv6W70ABGYOwQ8ULUNuN7nliS7Rw/z2
XDRNMAALUnDPCE8SkUxtgN8XQPBkuTlMPy2u18L5K6RuN3sbmyoeFZkQsyeqgBoS
6pG5W9wLySc3Nclmd8ns2xSvdQk1whV5ai5oQNLOb0g+fJmYlv6dHjOkh+Xf4qFl
e/Kk25wUjYYXbWjVT3eoIts3iQ+r4QdCSEN+h133vbII8FrdZkqcR5jgRS0c9wIx
mjaesIfYsf8WdCwVqNXM/OJApjcij3Y1kUMuPpadycbefDd82tmhaUxYnMNg/0k9
8g517mkTMBwuVLnj+neqVZNbcCRQ9Ocr3PHNMoDvfGmzKlqUTNrbvA3nBG8phzng
1oZtXOsRlp3MkiWe7M0At0j7mkOXER1dDDawRVdAQd++zzeUOgYc6eCrodKlPvg8
6iJvsj4+Y4WgaNDqcnr271W3jiSL7jEOXgMzVYPN7EbTDh5toA+9Dd05qUtw7wxE
OsB62q/hNyezl1P5xpA9qkMDnjWZk0l7Q8PwK5NwLES5tr1o1Nn4nBsDo8+GoJGl
9/HvWsqz6wJA7Nak3LzS8P5n8Aukuxn5H+WqaUMLLRT3BZwuUjRdtbf/nTKyA5Bl
ERDZzxTs+4J1/Q2EPJSJNhLvnteAQORBlPaZUphdWkv4Gcd0DqpM1AdOtzFcdh79
pvyd60nAI0XhNAqfjN/tasjlPEVXerb+gMYu53VZc0QF79OtJL96uFnAoXOL7tgE
ruvVXxOwraP1uPNh6jUBditj7FlmughE9px7e+AhWNdMIin7ZK0HdM6938Yy5gMb
n13wbaWLlZSUl9SRstCyMl4A2O4DXKDKeVyPL2be6QR70kMnODID2nFo1ixZF6gK
l0r4WgSugLBJz+22xPexP7o/arQGmDSWThTrF5AVQycoRvjyDH0Yzgkl3ym6jHNy
jYEOZM+vHIr1EbIj1EWYXS7cXq6fcBGUQGMh6DeDofSvEw/C0hDJU+yby4JP7QjW
QSXh2BSzpboDvvOgk2l/Fmco/POQO5LkRjwbdFO5iQ4Y3mHGVXM/unmwYxHpLDnu
MBzQOhIZTFRtyAoBA8mD+YJDjUW4yPA1OLoLBo1umlm6iNwSx64XDm12mkaLc+Aq
mQjvwUm9Fuvx63DvXsXsMGQCzoc0OeUkbzxgVqqb08B0WoUj0CUKT4PrUKIuYHQj
XzOPqRb1HZi/RD6GMiSs8/Ctd8cKa3GGZaL17Pu1hEfcRKx+8yQ6MxVQchzY6Qsv
Yh/RiXhtuCwzn+mCUoxcqTnvds7Y/DqMPOFssYkPq3HQ2wyqdMvt/Ctl/dm5l+t0
OwRZojep6qiN3uaazgkox6hPJ7SnIRstg1VYbixY10nrj3eexKX2w99FIeR8Y9Lw
O4OpsJGIIeJU1u22TUJ/c64IK8MnoiWKAPmRtQfjWZUt6ix71RadePs98v/cXMFZ
ji8szsfBaiTxQyZRlQ9ZQhnRxOVVRP+qoshGMtnml+jffaAmervZ6rL1pcKfiY34
cUkF9fUO0aXo6snk6Q9s5Tac0fjiJnX0EbP5OAm1IRCFEy8RMjjX8rba7bduk2mD
rJyQts9f22Trg7Wk3/I7CtHHzk61PcfZMc/Kbtm28AhYZ0BDWYqws++1nz3iRKGS
p7DA1dc2xD63o4cytWVo3p3cHOAcUdPomS9CYHcyZ26Di5OaGL7H5fQ7BReESb6X
eq0eHABwAhrNbMYx988pzfRB88Gb4wAgTzf5r4o6mMRd/9RPVYFbf8SNqXE7PYi+
RNlwpAK/PnemkC7JNv3FoM/bBvdl0qYZ56G6E4FFKcLuH5WEMDe+AqqAafinOncR
hAqX543jD5zob/fQtrOpd2Bxbs5IDbM86HBUmR4WW/BDpKO1EikvZSwYR9+J7hBe
cCBnYJaDkZd0fyG0Sq+g6fMgk4qklhrxqlbhXHzhQGwIKf7SsbaDFYohKPa86YVS
DcWmh6W2S2JDy35+pym7tQBh39Up0uCP7lYKzc6aNIP4EGomvjUt4HJSag5aOWMg
N+qbU3l5dv/58/5JPqrHLpw95/iZqAqVJGXb9HEc72r36bLcKM+DVl1lw6PymUs4
3bKFSgPSR8aDoT+RV4Wq0RUhHeXlgkuwj5H6MOhXhI8t8K8DSumBLGTWSWnskLbX
UvvzmZvpAIwmux2QmrH2QlbUWTb2Fdc5gIna0zDRISzhKO+Fyin7BhsEUlVmjFjT
2p2PTSeGy1/ddyVteHRy21KaQ+S5G8pqZW1KBvLM3ZaWdlH3a7LIWg8JDTnoKhcB
E1miTDj/B3aey/NMuqk714/YJSyU8IibnQ7Erx2ywjLmnen4zK5M+rFY0r8qdy3s
7grRRDZZfY98Kcz8e2hPx6kzGF74g6/zV7VlU7mtlHw37Y5PMEXsPGNIyX2yXXbz
qhv1O9c94Q5NqqbmrZRPjsVz1An9C/fjrzLbOP0+tBojiEOy+Xqp5ebRhc5budZ4
lUM7nEtk7L5Ejv/+H40448Sf3VbSQmf+Tz6oooJQkYE1KJxW3uw/E2GhJnI4WHdh
W0YNJnVx351rfzOrUcIMe5paVWSMaRC2pE7niS5GSui0pm/v2SIMFi73K5VKJ68I
BF+aoGsCL9gN0QH22irTr4D1F3aYpTU6tGR2PmVnnZjJvgGdJGToh1Vd40QeckbI
PAKu+SKJLIGmXrlRJ2qwDt35MduOgwgGtfrrWF+4G6sobgmJOR/D6w3s3ihBezsb
uejia0YEKltXn8jJ1lRmsXakSzghKKX04OjEBtCqy/2EYRE6HPveQdLhyXMrZlTp
tGEAQexv6roXKyHgyc6mPPKsm3NlFPvU4f+pBEYVpgRvrR8g3tztf9nrzNcT582j
Uec97ulPy/yWkKoddHmKNntjfrqdInJOyMAZLddSIGWiKspMdCK13PGrFUACqrgb
YaMEBYbtWs65ovtJs36zP+Xm/eS3M0k/KdNViAR7LYb4DyGtSm3nYGnfBypXy1iB
ZUgYam3whA4UvjHRiA8gQmlit96+mjBh4pd/g9u/QYGbpfKrYu7ld+WtDwVu5N/K
xFlod1aEqjJnxo+neHbK3YrVFSekT4Y2sw4BEu9fXAx5u4LUHhobjruRbHji2OBk
bQjbLP8tmG6VJQQKvwdI7NMinP00jYYx30DC58wTsZvR2KE6A77Am0Fvj6bsiiaZ
kUPXze3LuD5al4q/6/+4kHf7dA71ymZrpC+zMLvEQv/u/ZYv9gOkNLOpvyh5Gl2y
3osTWtRZTtv2wm9dRhV/CO2auslmu9B4y+Nb0k0vq/wrpPXYBmN0W1IMA4V9gZej
z1t4TLvCGRHQ7qrsc+pe+tDvES3amNCx7F/oWr9ZbWcKU3c7jtb/80+VsKJ791Cr
djAuw79okrmbNCuzWd2U6w5yOaJta91/Z8pJmLfi4Zb1vlC1mRV3P2hva9bo/6jJ
BWbLt+WzL8JcrEyIrmS8b07HFese2ajqaEbKNAlfSvDyRjLJhB3a6ubarMchg69i
qm0dCndrwkKdiYjokEiQV4uLgz9wGOOx4fdqThU5DUEPFkVN0qVesg46cylEKNLg
H0Qgb/NKZPbBqYlY45wA+L7ymNLHMx8oGlXDWM9W8qqcotk1bI3Q9LozcxqnVKug
VNyk7NehYcayuZmi8XDdN7rJgNdf3Mk/lcE9BrCvGUqLFgQcoWLvJYlB1sl4iebN
UBQlMgdDrNiko55VBEKsP6svMESm/CN8UTC84E19IRvX/tm+eioghNSnPNOUMzdF
SwVegLh5lifVMNS/zO5soycyPGJIGK/w4+L9g9BDeSScK1Xn1vaGY1fqdGOHf4H8
qwYXKehSfyCIKiDt+5RqW1k6lT2Tvmth8UGQc9xh0mWmktBrUmZv+F3H79xe4k4d
JSo6UAygQOFKhptaBI1Hdp/N2vZCVrw9sEj8Ru0tWLkIA9v+s62MzkXent4iIcqQ
M6s9/QMm9YjTmz2ZLTzlWphv9T95D2BAEZL3Hdj9UkVGtmCNLsf3yrVToBKMBtXl
heGxy8nOQVWO6LJMNPM4ImIbwAv+q3rJNlBe8Stop2oKQO1CeCStW8w3HOzVodwe
G7+r4wfiTnfmj4a7SPOttq/DAV8tjJMFFM+pbY/52gM1Omy955JaPf4P2OftLb/t
gp1jhU3+OTKKWh8Fkd+GJ7o9uvFxZ4sb8wjHwdVOAKn98z6uq+d3lttFtC592ml9
h5jqtPw61nmnrD3ePGQnSK8p0CyfmtTJkRIW4pj0C3FEBB4sfRZf2qP6juSdQGjj
AwEB2qctECPmarz3BH1gmSw4V4Bc0qYFCbb747iQZsUbXwlizJxLoBZBCUnhJBwA
NAQZL+Kcvxmev0QQXYKk+m3hYkKl5VFkHMw+AvWKKi8fdv2WxGQfeZIK0/b5ZMfO
zlXA+OkRQuvNVehPOyDEwu8P5WqV6c+kus9DlDCl/ZiWVGMNxg2MiuM33Ca1yhSI
mGa0rx3q8jtIdZfqB6mHjszZAw9tmGhBUvjKwo0M0IzWclr4ZZUu8axFgR2tRgSA
q/acH1vqglBKneqBBrbQvGTtuQSuv0s+AXuQWbcoB1cXCe9G1KmP+sON6Eaoir2D
/XCJQi3EeVXGg66BmloFFeFVKLqmfUZ1C5nNDK+77p+QGTcfvg3lHKa1lCHctDYG
S40pKjA1Nw8nR23iif6EuEvSnFZwT53aIl/9HSADm+JH31riaMqOow6a9O6KNiuP
ytEAcFm+W6EMFKvYva2lnenNu2TCx/Xho3q9eHOpRW2nzk2uCZwY/b91gGmP2zHW
3/m1r9Q7TGf9kDMhPGrysg2pmvjBf8u+IjjA/iXXQlP+rMgpBJ/0Uj3ABJHTWjvI
I2d/4bkMc2hQ0jYfSnUd/0SNQSip/esTo9g8cu3I6zJNuIibDiv/9/5gbZ3D65kE
OoLje7Y4vfDIrvPI+BsBsZpmXv52e12uJejd56+kQLrcF+eRwk4itq/wX9z+rh3Z
lwX09pHrYV+FVsnjPmKyDqvVh8R+SUHTaQmTe533rEhNUeFt7wgswN51Q5yoGZjP
OXvTsR+rhHpW/9jTunr7HU9wcFgez/qhPYkaem3qhd4GaLgdD8qcb/s5pWgOAOHc
eNAKVwUAVQ0qALz1ehC0a7R6kqbP40rMv5d0WF4fbsSebpP/BD9bbtJ1fP4oT1lz
plxFN6IOw5DFdpkeny+1/qpRIOI75NRPkOELnar4Nprr0WlaCGhA5MWv8nZ/cx0Q
77mN+JlQQL7Wq9UL/Ct0ZjFrIPkQ2BFkUTDGcwrs6eZM2yobaj2X1/Fc5Dpwv09l
zTNmXZrVMk+USc07srnCQiTctJ8FujRthAiB6SI6Vjga2vdvRJ97IG6jh0Jp+Kjk
fMY3+wXnJe7iyfNXmKM+jx8Wc2kOikdOfL2NwxjpSJSPs/YetB9XWIjqbYHqBMyj
42Gv0pNsKR9GuogIerQGd+v0CZxpMLe1pktNSDKoSDVA0MoUYN42KJmDmt0LB8X3
Tt30+OpvJFUH4xgGrrf2yUKld/kmciX5glh120B0GCbfpKHpEo1JZMUYxLN+94vu
QCbdA58CECvmd3iIVdqGcm2WchesP5qOBVpG3cERupGhKDytXqCxI8kShb7Z+d+l
/25KzNMfm3KE+RzHt80wxt5t+7n/BqJSlMNwzvQs8jPZSCO9bBhW5cR/EqJIcv5w
WRIzAb8gMXCPJc6JrGT36lDRERIK1rxRDog+O5t7siUJG7paD9fHAlvs4Q1squOk
PVlezwu5XsMLDAKvZIhrnpbRwJuPxPaBUDe8gV6kenDsy6dM+iO8V0ujkTK0xwaJ
6kFS7XTW/A6FkMJpxeeOQoAEX9vnmJmL9o99gtK45N3/A368QkdamhBMYdSUknci
U/qG/CVa66RTU47/xgO0rhXwARtkpv2Z6yR4O9nlQI3Qtb4z7T+Wvyy1ZLEY+9vO
hG+w7IIEI6i+o1aL69MJEbpDlTZI74MrmQ50Pkgf3WSnYNup2UwFErv38d8QLSw9
sCtgwKemcR3/HjwmMQW2SYBXUlTnJp0KkQg8+K72xuc37hNYOrWG5fp9gJZWQn++
gaNkt2ZLpf1mpGhjYNHedJ70eiDSbtekmfhiAaUt/Y+zalbT8kxyT4oze9KWycrD
tVIQw7AgvaLO647D9fiJToWVIorDittrRZF98QsBBkAqfRkYEyQS75mX8OqBrPL+
eWWLj1iojU7Y0Jw5Opde7/aIWNIghl5ACh0aGpeHJBSWC7yVZnYiqlIZS7HQN45S
2YndYSN1fG9cyuZ5COfTi/nsWD6rLVCK1qkMZzlGCiJoMx82LdhgqjTK/l1uTQ/y
BMgk24iAjwCefIpK8MKq6TJ9znGtIKr7xVZYaN4nW2lyMH+1To22g/HNNYPYcYkG
zPgObCh5+pCqxLdx0JtgU8WVoGU4K4JYVSko2zAbrceV02T7JgbwE/bFMEAtKLqb
NA4dCKaTKOTzOqUsnBaCQ19l8IzT0Ot9QNRSGtZirP6crxkQg+H3lsigFbJhLkdR
B6w77jJZ3/nwZ2gi9bEN+1aGMQ3UnNci9vFxhgEfMJXS37lgYg8W4TQ5UhBdLWYk
lqTMM2W6NZdtB9JWiPm1MaG4lS6V/WQw0uge1NLIqGHUK/LIidlZzo9IO+VsPyPE
e2p04FFHYvJqC0CTwnztUcHO6YUKqMxKyvvKw+WBSxbx6Dmp9vp7vx7opvaY6G3A
oCMrJeknZU9EV7suQd3rNRLf+6mi1JdIONlHjzpgPjoc5PNvkGB7KMSYLU1opBRK
nDxs4y8oOupDMAehUD8W3qRnuumB4tDU5V+LZU3k6s2now3s2e86wlE3axM/IOIT
Ah/RiVHtginZGu6eC83x6LX10lnyYiZzs9hpBSAvnUcV4/M5wVDnABbmZL/2cRPj
32h5+a2P3QgvriOLQLhde8jvQYPuS7uWwjHQiGjorzhmhebZ1EBGHGU/MS7E6lFi
fks9RLYEm75waCn9x0gzlzr6ejOoluH8/8svIf9JEdC6AqscPU/nvZTYsjmo0xYt
QL/jsh1IEbHZw36xioZzNAB0bZFZEjz6IdMDbLEx9ORpGkW/w021bbJoHLebSana
PsSq7uH+tm3sgUfVDNFf3taMP1MQvuORLe5BEqLi3wShsBkADOPEe1dcuelf4Vt+
xRi0FqhjIpIP8FOvhctWX+e8Cl3mzF2ftvKYOWRubyS634gCc8Y11OscKHNE1OL+
8uGVK9IqHEfPbnA33Rcuag9/fMxXqoVTEjc3fcoLPFYfR7qcQZ8ZYMMq4wCBute6
/dcp6xaArbLlzSA1lbEL5dAQieAW9XMPdEJSyLE7ckIiYp8VTMP9m1gNktWect4w
+BcOtysAz5C43x3ZVJkjXdaJl0fylufxwOX2oI1He6aPMhXPxtvLR2nFCLPbOIND
WziWbkeknbYfTnpAVzfCNIoji2nGjkEe7qnn4ZWdhhtiUgzjiAYBQ+WvpiLWF9QL
oz+FwxlwzHkrbN3zEsiEMDiXI4lQz6GeHEyvz8gmD0k788wU7E/B9n3Z5nkSHuoa
Y301Q7ArRIi1INsJiSpPaRfMOnMEAeO7OMH8v51Mo7gCnDXAuVNLZ2pQqlA99AUt
1PQjCt4zGRa67jXr6BC0YdNQFHmoHif/ohEkHhRpX9I6szBrVFqTqNKgU9vAJUgi
Cuv+2Y0G9OC951/vOll10z4e296u1uBaE5wCe3wuoV3Eem7TNYWuZx6+rwduvEOm
l/Doand4Uit8ap/reWFfrzE61A+iD1ese08ON0brZz4oTtRHcD+Q3xa5i6q09nTJ
wB2LRtyk4Gj2eL30aQ3nE15tM3jHw1LPDN9l0P0Rll3rYsGgrEO0c/NpaFrVlYQi
5BTZ3lRMYBA3NMhEndhhy+I0P9PqzErU0kxauG9yKG/17L1ThWIpRN/f2eQ2Rw1P
141MHpKRSPUSGOoCXz646Xvo/Kc663EkaYFv59ZHkLiIaWxnnLrio6qN4onRsY97
1YZ1KDW1m6AwmZPYuXULIydTyib/IowpAYgMOuFeCTScLjKcIOS+PQYa/TCzZTqf
M8/MAwSd5AEJuqtak0e5pakx4iQbIMBEH4+9z9S6tQV8z8WkkI7StAc+ev9a8SJp
i3DUDPO/vz8YCn8emc9FynXMko/p5AG1lOJtb6uCppQ2NKNjJTrzcKsTqxZmQLg6
C0v7HboIICl8STiWvKYm4H3ekpiJSkFBls/VomLbLDKyJKswwgb5Pj4OrCyZgSha
4dMgPGU5baZbNVTk94SJ//dXBp4AD7tubdM6rRfCePbhSs99CO1EZLRYWWhR6/sV
RMSmdb7ObY4BiQ7DzUV5hao7EGGzHwQsr7QZpqf68frFO3AWHRtT4+LZEtoak6nh
oePdB2admrgarlfP2ls7ydn2ik1pY35dkkMoavl1vc1gFHC57G35hu2fW33F16tW
691YxYv4eOZOdDhqQ49/JFuYzIera8dNAG/spkw3lLiwMx3PEYHlT5gEyfIb0zO+
NWzLNx3gGSdEwmajGZ3XRcJPoMB5k2BtHdKYErS7Yf4BnBb/aIvk73/WoC7ynofp
46waRefBEp1Hi41J70S3eVg3yaB9rlDF9KwdYJjazDtN+TqtoyqLVrKgiNZwFuTW
YtcxAZPQUhJKYFrVjE+gLVT/6eGNJkxikuN59QS+sfr1qsDvq3dbrFtbiqzaDQtJ
zhGAhl1v71cPjLdkdruRHBOctlAgAscuvBxSlXhP2VvRN00uXl5YKeWYHjWTO04w
c21IejS3UTxoSoKV/lOqJYM8ixYXQfAy1TWn3LlS/0yyWOr9H7InnboC0J0olGt0
AJBfbiwwdsy6y42X41FK2LqUOazpJVil6QmgRAwFRFRp/W0u7q/mrvo+ZKFt3Z7O
rjtlx7oULVB4XrJNc1pBPkWybcym/ZFUfAAhwIWilrcqQwozKyeQdWBpv2hRlp0p
izA40YW2l8g9IiPWOZzz5vu7oWyDh4vJxaBqaL1Xxd5iBIR+7HS3n1IbR34onxF5
Sc4x/oRLyzv70BMXCZZKCLZqyMFn4y27TebeRpoyyRdcBpDsuJvLnyNsikUypErq
xuFyJ4zFq1zzN9esK//jOOPMf6lkO38PzLQWKJZ/xDEHs28mU9mCk92EVDEtiKW9
sQ7DKsMtzO9S70yUXWwQABk2F74ZBBCLCw2IHnO2ZUxblRtG/vIEbSICarPpkjG6
UT2BhKprqnrCg3KxfEJLj3DyGj3V+7g10UFm23C1u3qICn2p1FtQzq//su9ylumb
bgaHVayFrVgSXxAHOcd9AGFFZp5sLnp/GyIasBZ218EGQCOUwDHKzb2lVARbcxqu
9Zj16fi9Gj/wCsOyyn6cbgbTPgVesoKAsPJC/Xm6ETaWPPnOkV+8sQBG/rB3kZ1v
BOQy/dT70tuvYVd/g2af84+OzbBzA/a80rsoRPTY0jBjBSfX2FRRDdVBPE+rQdHV
BSkcThIdU5pUPAGTwwPFBbbbX3EKtjKJD09fvO4aNMRQGpEpLl/H5gYnz6gpku3R
fLs1mGQ5uAOGdc6BkV9/d0DnUExCNKPX57ovQdWlM5ueZGHfXq3RWIFKMJd8uiBQ
UFBG9dIy9ozkZV58mrYphF5lYemaWPVtLD8wfh5HGYPB4uh1DlijkrcTBurvdgxO
P0FbD7aHsXj6yNKg0qSDhDFLoYEKVeBVQ9GF7dxg6o6YznM+Ts4Ale681s9nb0cK
OYY68vkpgeD9SIGTW65F+hzrOSe6HyhVD5rHE8qTPUo8xIcFDbOqZl/NSLkdpsL0
kPQBKa6UWbgVwwX0OK0CbxmUhCTgFW6ybGj6yXguehR8gRv6NnMWvZwxRV6PvSLW
Pkck+wj2qswFxaiTBTeZPuu/LTIaQm3FsnpSowsSdyQjinvM3y/rJ0zzcSqqTpo2
2BekG+mBwxQBPyT5hzUllPvR5L5jOvS7xzg0PcA5YwEokx0qHFLoMuP9kvq3qelf
ILdCdU3wFpQ+JdkTq0nlePFQqtaJD8yMalwAKdLodHTUsNxrCeFfO2SIfvnaBhl7
E/xQubDO/HZ70lFo6c+7d4Um3uUaY9Kmjddoky8/8QdUiOGco6Cd+wC5zqrMNPR2
nnrw5tvflnaw5n1hz9vIm5V2p05lIPv2EwUGMTeV7/4AwHhcEO/HXBC4q5yGau9p
4oZdSswe/Bd6gWk4N46DQEAl/upMYdmdTkmAocnOhhPNvxcQD/l4LyipcsTEsU8W
wt2p6b0bSTKmCstdURM7Qh34speCNJa4Cu2kJDVJdF7u1HIOBcdXqC8YnZTpbcr2
Va9VSfJ+jyTtmd2aD37Anr0iwaoWE4sZDtLG11jrr4xiJrNHxTL5FFpLPaSkqX83
1Ex8ic/n6B/aqj3y1I7IiN/hPUTrRZTT2r9Vo+GZ+n+Amklcq505xBa7Tx9DlkFV
5tSO/srp0DyBlmcOGQG6TVWAxPfnQoughvCyQ0guR4Aysbg0KWzlEUdOWMVmUhSx
WEr1ggrjXlyyjjRc1iZJNzCB7unsg09yhYEepDV56tLXWNenDhY1hD21LzJ8iS52
DWJXEnuguzejCzwrJvkO59vRRqSd2QG+FJWrPmD1JVZLfuPsqMcIKDoDM1GnsYD0
Dkss8g2p1U2NUSBIOeOteNtf36GeuANeRQuHGrpq0MX4YpjBQ2ZOeqiYFYtBVVV3
6dYs0AmQVHjHm4UNQ56FXgKiweKY6rvt2FMiMV9ZGg6J842v4sR4qrZ1Q4WFd/uh
Z5gojzxTv9OHDRs4LT97kwv+CXHVh+9ub+yPnNyww+EyJERkiQqp9DG+YfJO5mKR
On7VdELS6HXvA+EF9Zd3mi83XQPOTzuXV0YMHAdPYT3JBKwNDmc/D3U/puxw2xYK
Yyq1uChdlTUOC8wSw8hr2UyNQ64xOTKv0TLsyjmuBkFsub99YgBGGf04NOU00sTZ
6vkrMHbfOOvoSuduRNhxMLf3u6cGkUto96DeOn1o3KNkJRwd2eXlFLn+0GsaLoXs
u80zmVZbGzYfjPtkrPCXCqFxezfB+ewNea/FXB/5pU4v28zmmILs8/e3FXQP6B09
o/GHU/VIUJm6Dojwc5jZ299Mqp+6gL/QBJhVlTBueWld6pbSqhmS3exXa9HKzxyW
vq+as1nppq3X4O600/P9wh5HeBb+2/d+WCThN6dnr5gm8tY+ha53W8dPzUjuGFGi
w4uA0kNhTLxEK4JTLBQkj9K3c7OcpIRTGJ7OGgo2j0af2F74E2Gh5AYr7wtWteDH
WRwyrqTwtPAVofaZwaBUlki00bRCymTjOA+BOL7rrI8I9EqsAVVcyKV8kPFhXK0o
lFoUzlACdXags861QsQRN8u79HaLqs7mG8FSdTDQxBcNraYqmMPsHFRfyN7eB7wz
yHaVN7RgbA+sxa7tsftdWGvQjl9wGUeQ5cmOdUZ6HKmx4xrNyjncC5H1QJ3Mm0vv
u4aXmOTUmkQvUPtLzo1G0g/2hxjRKq2QUDaidjR4KOHCOse66cPxN+0wlWkLGSmI
0XK9H//Nob7xZOMhieg18DNxvnR87jwyjPcg9n0GyjGeXBtkzviB2nBLmarv/0F5
F/FC4Sl1odmBzCr8B5Flvd3JIRnopB4H0mBBX5P/87Nq5lZSX0QBFqYuCe4P6z7i
z3fgEzpAYkfdRdDytHoY0fFQzsaTs20UekgGMKbaTCnrWGfGWo8DLTLye8/eaVB0
phrkv+ShckE9QCKJhqEVUKO7BctXDKR/BbKwXE/w0gdpAtFeYBfHwees2jnfLofJ
/42mvXPWLsdsj5aWvIeoCUrQcZGO8nQM2nIAbrP8QeElTOghLzxyXcU9ZyQ9/Nu0
6oPFh81S2+FQgKi+kn41YzUpPDNQ4w19r59H04uJ5PBlcNxJDe2QaPVIP0exbv9c
q4QImbFDFN+2vM2QRTj6EHvN3IQF+wlf3rCNwASxu149zh98FyfgSQjTU7DGkpTq
2lr7DnkKSUZD7FktwtSmnKPlGDhKz1/PeCNDgY4z3AbEJ68xHPuxHfduIpPJMKpZ
4pkgOAZZrdCnJMsZ+8z/KlOVlXDliSEo+jlcFV1I7tH99nsF1ZpXseQud8l6Qn5K
bxm/V65OzjUN8GLoqkpH/ifVqmnZCjd85FqlCDkGxih25ofmJaRwn4FUCPtqPCNa
XGnOyxKJVIDXkFShkiJtuJQUgsvJq0njkhU5QsnNDOqn8k3ER/imHaSkc17HCBVX
hQJWwGpo1aH+lkDBbjV/kxMIZdgkWGiEdMAizmowEBn+qJ7KjNFSTu41fg2d/7WA
2nhwcb+mplEE47f5GtDc3ohSPVZm233OPRV3298YcQLOuDl7GDg1Y1hPeDhOE0kQ
nOHnA2scAe8YJZzgAxm2S3WRN+r5oh8rxlNYwBX95Z3a9Pdp80p08R/JJqunUS/y
IaHjGN39nPrIDaCUhfkoG6KUVU6TqXNyvn6tchSaV8DBjfLGWTtJS24E+ghALROW
FozJq6nNztrYBSfhWecBCK97dxOWAtk5K6M+k2uB5fguQWc/ROWG18WfymFo+0z0
oycpYD+G4sI7UOs6PNMaDqT/CbCHDCAsrV1SkFKDkNFi6gyDzilxe/lx5iJ+HBdH
iEq+rp8pNwNYmgOCg9vqY/smur4BVG9PAbF2bizsO7E/aTjyKMSB7kPHko0yqJRv
AQVe+O6+5wg/bb8UN8Nt/MhjmnGlf3QdWROBTZlQ9qAMRtrH460XH8iqLr5LI9Ih
vDYavYhtAjPqpNmtVyaoyU9Z9bj9PmFEPgL3nGIjxN7T1ym3Q+Qv6tOaIv/LwgPc
o3MW41+1o8tZXayxHiDLRPQpy0P42SAfNStXqAwaMuxFbY1ihFlJCAfhMsIHF/C+
VblR5+5VXFVXZeUIwyqnOyG2DgPve0OajCfMQ+rJFG/OJby8d+Q8CqeKhJe3G1wG
FbbD0W+59RMB7vpDopV6KH0B8Cbt/Ne+5H9oFB8o+ZbhoxI3ssupPNvv3zWV+oJR
X18Sb67TkNaBcoOph44iAifKuFD7Rfbu4ky339lB5kyBwonIH2s5QhIIJA+xbnFV
uG0MUWGliAN25nlUOCs3j9UvJSJHcHKVdbrA2sa822QFutiD6v1dWWkvhlkddEel
BxAnJx9YS0S0hRBiitJLxnmJuLuR2DjuDpHAcKIOlDDZseHt4tbLlj33nJV2JhV7
gPXL9XJi8ZXJTajgFRNbOykBZBjJTwFF+8O6FiufXUj+alS/R3M1hekXr6X1OUyb
bQby2SpOKrmySjphNVmz7nK5dYP3+2ZP/aVExsmiwBrDLANBMMFom7f9tV4qOyoD
J/zamoXqDWq9KfcAFjI5j1c3jF9ZUgWPC0usYmxBVHhuHB3uIwI5LubZazI/PvMq
cjz01DhreudM9AXZW+N0ObN75ZhFQncfZQC+U8F/It8Wxw7wz4aN1+YflulFZyIv
GT1OBXCUSeXFL/guqC6jsF5ywQIxh5Fqsl6QVkr4i70LsjWhuf1yEmICgzKK1mZD
/2bH0BaO0GMdHQXg4ofUvApJ128HUrA10pLBowXpiKAZ+yxJ1BwQVxVsNFvw4FKa
sfyFJfuK055Y8/3+Z4Dzu5Fbr2Pxmii35KubUsPMOiu/MtckMCV9x/GD1uFwAf1M
+pzKT5yKW6x1wdrWJrwny9QYt6e3282ScdGlTiktqokwDGpXTtrPXpBehTNF82lp
ANLorZotkmr1dVD0nhZ/WSCHTwy6f7+ftYr299NNnkiX8CjuX5goQrcPnxVvNaig
k5ariVJLs3yMT9YHyEfFsBMDjaNVx8Wi6LEy3at985rpTqJU/UfJuovLFf7YZiWs
M/IRaIlQlRjJEE60SYhR8e5quRV+XM/3xOwnADrp4V6vWAHIDbovU6TqsEL4zAk6
oY9b7fAzKCcHRospmldunhK3lojNjlJD2bfWA9uTbK9NSOA701myPH2jQKLA1rif
AxBEFtLpP2KkPESCzwJcofh3NmtHVZTw75lfX0IGyolOwn+S6trPw74a0BzmLYd1
RY3ekc8WVezu94qGgjqSIp7raiVqw5hVRyyWAo45LOyGGznzkNG7CUS4C4JZpTQT
1mRnuX7I/ztPolxxlynBRUbEK8Yw99zNNdWqC9QLrlOQsJCpxR8bWjKR/30yjU/M
hx7v/bupbvuEchQyd9RN+v2TtMhmODSDHpPK99/OnHFMajoWauSa8f0vOKIHz7Ek
a9wA1gYYMhOSZz4XCC6Rel+++eYUQDxldMMIfcCPx0w5Jo1ZB/F2Rp5pPOckNq4K
FoxAzSJL5dFTXJizGHrLA3kwqxmCuFlNr2DaM2ejXmzOqkPzg4ktlxrhBgLKcGv9
sNa0pxQ2p2tuCdXq09y4GL/HwtcHKfXdTCnQybkW80A6nVrBkwHCZyGoPss9fG+y
tKuA41gZp1ZW4smUJAK7drMqe7WCcKGYm5T3fv31opuncI8cfBj5XVYkww+UyRZl
jRIbPQi8cUKdwcdDmmhwGVdYPDJ5KZPyRevr4rECwifUWurfYVrATcrN6OqVFeQ+
20whbzB+EMJ7XvYvU0kZNMPfgQ331w41Cc/sATIwoXQ/y+pk2d6N9wbqO885ejBw
r9TgTgXr0HDEUZXElceteFhQ9sCcvIowbbTtjgZBfwhL85+P1TCtCPXX64zu9Cvw
Az6PLFWJ7oitDeTv4LQVyM/0L8TLLh2EpEv35349JerGVotJb5+MvlxNkKLw/1C3
6rJ1JZkgEyrR8m8AE3DR0U+kkTrkD2r86DBOUQLzL0Z01jICvLRvmTI5q+QsgFjQ
rhP6sgYitFNwXMXca+Zq90RZBTtfzLjZP/Xs0YJvBSLghFChK+T1yAt7uwVCxGnE
b5KGpw2xcadm2yt99/yZyJbCaVBIlrOQUb4IJ7DOO03tik2M6LEjhPZVKmeGxWLL
9T0Koph4O3xs/PAHlPrq7cahSbq2Ogj3qAO7icAOEe0Y9SqRDxER5EKSilkqdUHg
tAxbzCq5+fYwcxG+3UXzZwyiV0N1Rb2mRyGF87h+mVdVF9mtRnb0qCgRYjhrwIGy
H69TpKVx82hNqLHVvm0+YUYPaAEUGHXVt59pqAbzknu9jy6Mpf8sbsQJVqgqANVm
AOf8ZOJTEpGc33XgH6XYuP5h8HTbQ/Ps7v9+8ID9g4ciiVz0tzjyFPglgROExIyn
w0czJbWjhcnDKWVp/7Q+BJQJTau31oTkOuJkhp9XgDxkHGe7fA3Ph9/t8Ypi2xF6
baFWlDrj9MJJXNrzKabbh/iffUexwsl2IHolwuRkAXEIoUnn79M4h3+21+T4jggt
i8GsG0ya/ASmrhy7q8nA+vY9iwNfzA4Rk4szyeuVnaDhXPJjoEh3Pf46SFnhmpHa
jpwxdJJZra5AjmSnSCPWhLvrTvKrQScyaetnKopypwIDbbWbq833NebWqmbgCmpL
6QocYSQZHNLRcDdJnTqQUWD2sIiQIkTaUs8VEjjbesYkU2bloy4+6RklfD8j1OJx
/NcWP+PVq/1qY2cVYUAy43UNzwf9i7rl/izGzt2we5YNSoxLGWp1C35zieQACz5W
I6Zw6Q8Wa/K7J5EjTwEsYE9G3eo/ifvttnT8PSDLeRGSqOgT0bGJvD/ADnoLJa97
FiH7eN2ugQtclfNlJXOZQI4o5F/6+Ajb5B+X8mlQdSoLAtfSg9pCNtqG6luGHXHA
IUf7oYLiZsZePvMPgPCocEBXwdoIcxfMLwfU9SjJO1bEK3Jxr4i2zI7GQRID83MV
eKlwPobunATmgBY7gh9r9NAExBP63oXb7sHBczrOnWJ72sxl31DCK9A07vmytSYB
rgiHqZRJdSc0UypNUv7qucPAB9H6grEsfbZA/xkFsuNrYK6Hzk4bbEK2ccyUfxxj
3vIZ/Lm8NHq4Hs9VKLzptwfAQNUgkEd9duRtoLonYLuZ2ASnkG2+PBTPAHRR3Q4r
zXTXobrBPXvgH/39kw5rZlZjOHvRAgCb8rmKEcuoJgjPvL1HdHtCrKsQC/d5iLsC
duaBbV9BFoLwzb8uHAYbzi0ZDYVrcMifdt/w4v2BWLaxjH/7n3RCUfNisE7Qv5cS
9bdiUxyCNhDhlxSPJZE6uZWoY2v0+CTOBXbGC2O133vImZ1LNtexKR1KABErr6E2
rvh1y+/R4nXKLAtsOu2lszuOoQMCzYlj3ASXJ+3V0aYLU2mmrbQaOBN6Yvot6K/6
MtAXETLAMgCHS8js3wOEvL49RRdbU5CcEmw9LdvDPJHN1icjgpiIxc/diEOlwVSH
F9j9qnociyl+BQ3UDsjM4eNh/oEWgFffk0c2MyP+jRkaXO+RDV/qfDPoP9RZWUJm
FPCX2U6AnMYd3xr5yo+PpFo7uge6gp+kGNvDiEgjxGBJoENhM9EWw7UjOXGwwexN
2RwrR/Prwdp0V1yTeg5CxgRM4+NGHCDNAmb0Ii4rnUd8LtpEVc5bLiZ+WxL8qWjO
vq/uu6hiM28IrZ6cPZ2qq435KzMVgjEUjpn/mxtK9Ky1kV/ihlt+2Wqfz1ymkgW6
SFEoDPm42bRgZI7ognVHdTimjuSNF/QYK0STZgLpP7Zn2apb7adzk+/CzXk3r4nS
MON1KPuB5ZuOK9ZQcXBKAi1s5XlrW9A6ftCnNfj47ONFGBgvFpDl8BK5UgMvasfR
CWim1n/jBb6EEAvfaNedOtIHjNPV52BULEJo0iV0MzJnDpTTLWl3ju21TfdAuq8s
CfZq4OaKr7cTOtxebSIPe+GB70DFKl1CNdhFK8ofGo5IgQV+UKtm00vkf5Qckx7O
PmD1D9PpVvgUxbVtsaguGyVw3CSGG9E7D3WlqFuQNIBW+gLJ6+T+yAsGbzopS7LA
53XfZQwGkwkZENo9uUQyDFTL8iVwQy7s9alD4Lo4bZupD4s3Cc8sCV7tSe/kiziW
EqUcCdYrpysgvCi7wLG1IsTtGrIpQWzAPaHstgWMttBPQGnWfxnFchMRTUbdf26S
2I5zhh+Y1A7eBnIHyhdxOzmlNRE1Houues30lnZnaWu387vxZ5ZRbgyAOR5CgWQw
ZFSXys2nBwjc0sZHA1sG/6G+cRtkoklrHkB9+IFKKxujir7d9I4upTar9CZn9YPv
wT8/yDr4oEI6+EqULkjzTmWTv9yWt6hn1NjUlZ5VKBz1sbUd6zfjts69t34KXifE
12woSwq8csXuha4Km1KNSImb92rtxtQKtcK4Q807lCrPGsearvORVYaTSARF1aCT
tTrwE/sLOTI82o22LooIPQx4WjiTqTTZdB+5SNxz3OzAwDa9+ZzK4gb2BzpmgcI3
OJq5teAZaQhvg3klLxtGZ6SZ7T4ungAO3X5TPNd7MBdoUV0Ip2sAUnZoAnJxbUr8
smjhSdrZmvZBQD7oNfZKdU02dn7/PaLuz7BBnmfVGWE88ATR+cmUv4M2LFeTcm+T
7ZYdPYWsUYEdSX45ft/ri5/W6Y3gmHrLWi9P9OkEA5BNMtGg0qxkHuK3M6Mkg6KI
mxJgotdfqFRPQPKbboxlu4kP+YRH2b2IYqB3gpf78RXU1eMHGB4X/HwsjdxDorLl
H0974sqsFS9TDke18jMS05ct+l+6p77ZYbcfC6c1n2c2oh/aZ1RtiZ+Oi1pAjT/P
vq7ya/YM97ohR6nppuHXKizN8BjNB94Ji9MDSQhhfF+/5q7TL4dsiG2n4XR34tIg
dQDF2MQCk9gw3YVR9yveBv1LXcnPelNrNFHckIQ5Q3egY45ZZHrIQqhlxApk1QEB
3wwzOBkkbLPoUFt1gXk0ASaMkEIG4kY6wxNeVwdwMhip99wyoTfIyWNSkPKM6FTK
q1vOjpVoXlfY3PJritY3SgqiZJr1/iougzZs3YwKZR0EsIgYVz5PsDS9UtDkOVJA
4gT4t4D6JoMsA/qrnZeAJiyasLZHrNrUBHqaaJIfstlrysugpkZ3GmqJHKDfLsfu
1FsGOwfY/a5/tIh4I21T23sJv+b/AuHagpfYpiFOZr0JQ4/uwgzuOhAu2yQFp316
4uKp73fplen3p6Zlm4aC30RK3R145OIIdbSGLvAKhTxMokOEMTwyNH8MuIZ42ZDk
XHTOdqn9yMpSa/Bwp/BNNeuIc4NllzzYwtcV4HU9EFBxT2GHnd44IeRLXz6CZLCU
CEMniuhF4SWUohgpSDrjuIZWjqgR9QFnu0yiTgmj/sGVZzfawRbDhpsy6XURpBVb
gJcBUYF+hPN/pBtjrF1p5pX3lKJl2OWQtCusytt8/l/hH7o3/0kmKA1h7FE7lYm8
UEnAYb3JmNhmnW3QtyQzsdILAnOz3LJJBqzYjSiCeoBxJk3ZbtCVmJWGrYHTmKCr
37wVTbhCa48wjlQcFXris7zZ5ZXVvpmMMALoFvwNl2GnrbHlkbk5lzuo1BLKPeB8
Fvpj/jtzqV2aXPaQHRvPnIbAhU3UpcKHONu4JjNRYKJbTD8LybxlPoG0/ol4iw84
TZMD+iusIriyfGK1hWd/yDpzQ2JXjIOg9xcEtLxJSf12uLKQtw/I7NUabE80jGk/
c7aEzwRrNR6clUOu+XYVJ5mdxyrdtjyslnhuxGfoIP/vkV4yaLycenyE7PDCXEj8
W3RQCDXnazhGaQFQU1vAVduFrz3N+sfybLeSIYG4DzAUx+YiGIz2Y2nemGf93xzR
QAWCjEtgmyHsq6mxiWgr/l8pbTDGDz8UhEKnEaQot7asYHWnOGgpHyuNLOh42BHW
jIudPeq9jGXJKhJvc2ZnpCV/BpzD6snLdamaLs46JD+2kQWgT+iZ0yK/gVZT+vCF
oLvl+DjzN+LDo8hUUnc2F8y2u4vf/86fApO+fAXfc9pY6mOGwx0iZ8YXb/dqYKFb
PDniSDA30XD5Vu/ePAjUuQ1H6jdrcFSHqj6gqAE7u7GpKXPJJfR0ExxKCjHi42tg
cXUF1+bcedJEyYUMuvrWS/iRBKe7z0yoBiRJAeKnO4MU5+P54MMCT+/dG8jwZP3+
K8KZivLMunkMXXXn/uMXs0O+No6FJ0S9Z00kw8AlZHwj9gXLy1IUWHx0RPno3zHY
z8RGT1NNUk4WVTti7rcGDR+7HxpxogtL9tDtNDHP6rExS3BTw2s1lilZwNA+qTpy
EqHhkBL3+V6hCUZg1DRSQqIJxBLF+oMworen0erhYbYrQjoQ8l+Xzuzp5pQmhOek
NU+51I3qLVl9ervTwPRs2/hWmFFdhQWUtVS+aOPEl7QlfLVov9Alli6VIxV2P0ur
6J8rTCn99JxlJ5vMPqPLZur39nAXTXGCetBaY2Yc5MscNpXN7LSVoVWrCQwVbxTd
YwW5MbLz9/PHa7VCjW0VQgsGYSUYL8vXJ4hOt+VPEuPoN5QeqVrcgd3qRCr4nz9x
o5N4ZeZCyiePRTUEkxBsxNadny4Q5Wy9O611duqAcdaFaOqFaaqHp3WprxcIoQgk
YRTxdNuxK6BZayfbz1EAPhEo5wZKQ/5v0VjmffbYTWcKPLQEkZCaCA5hFH7D7yP+
8uzQKBcU0TjBLEpZHpxOuTkjiwVWBSv/85y1LjziORM/DbU3/Dy4+bFRQagqROJP
oVZMlUFnSOrR8B1adTLiFmpczUbUr6qg7MaKNwALmYQINp5EkL6jMEb+CM2SGz+T
hk9hHprldMumtxkCOQ517DgLVy3Gz6A+w3BBOoE0tDYsOh8Ga+98bVIff7t27iuQ
0WZUq5GrY8MTq9v2jVIMaPDGUhwnq0EbDqVW4zrzUNMQeDjhzvwpgNHbJYa/6C8H
Is7NmhJCMJWYmkpvdqIbm+jMlBhdGDy7DQknetcHXHT4oZpW8eiTUolFKnSkzQyS
sYsCFVpr0PLFA7it3ob88Jw7GRI85PMSxGVx9Y03l86IHfmXUthQrnKlBvUkhFOw
d87vPN8SB/HszhuaohBn7ZsOelEKau6qHdfQ6UL1TMEeIewjpYQwYofZqIfhmzHG
VJFzbcYEywKOadtGntYRDYMjXOafd8ptoIDSqLImwPSCGDWToPQC/t3LkNyMq70D
dI+lImcqmZ7AOXral7YjEqzJYZkz51COvWDlUAN36ZPUNjHciYBy8wcVoROgRxX2
MC70LaHQIbchv+l5PmQz2Ao1dZvzWBlSEmLZn0hKrsny6YtCtlLghzJr4DNIobCo
ehOu+LHyqSc6FGVkzzlYTBpYvdOdcQh+lN0+7rFis0C+TOT412u+3Ntthw5Gz3QU
lW5317plrmq4hSEvdRy0eF4s8pMfp2iYoJ9Op4Dj5O8SKNHCDcHoGCzukhvnb6zB
buh4frSX3iX6cBmh42jN9VvKB/rWu5xBF183gwXoFGXaXLRJNyJwp67fri9td4pe
nUnQc+QyRej6WKywg9RAynNuALrXQZv820QGcJfsdG8UEM1Hyim989wX50emKCwL
bNZuQtGXeXuzegChCVzV+nB9zjUocKWNBoTPMg28WBNK50uuS9bm6Pv5POw8oP4Y
vm0W1EeRjDT4iHEOd2Dg64zqLnmYyrYdtpJqsuZs8a1ZS6LtouKdMCux5MmVaSam
/n1gZLF6FtBf+XxDZ7GW36SiGAEUpFWFk/nyypzf4RXLsLuwjQqupPTY56AChh9A
3d15ZfoJT16fn8yqV/vmzrxGD8x2bnSmDxmCsUXDKo5RTd1YnKsPnRSJz0L/1nts
UBPJsx4SXIYWbpryWpJswJ/jvmfUF7qCDz0nyK4kQo8oD7CJwAx2B3T2JyjNa0kU
OZdIdjfqhbLwNjseEuHhN1935FWmyo4JrbLdWWmflY9NdpPJJIGV5JYltijYOV4v
dxrN6bXjVWF3wOfpGTjwpyphL8uWI833XFbALn8bwSfgx/UrDVjXvgqeuy89Ot3g
N+NGxhFvxBC+HhVo4WIQ+fPAzdS1O5VA8455iqVuAWVOv7J6L+9NtdwpTzB/TYBN
Hb+LvheDVa4tLwxrIB7W/1qoXeALaykBCzcAOeGvYDRZfbh54LujneIwD3Bx8qLK
0DNdMuWmKfeq5x+tY4m+0viRZDsBFEKE/jjROLSSVtbPyDA0XExlE1/qBw5hptdD
2jKHwDwmNn2qBtwx4xsEg4WoWarmWUlpe+6Hkz4EP8kQoTG7yR7i91ieoVnQhwLq
8JTRTQi3aPdcZQziATagIFGezo8xX2TGriKrLoA0jYDBOIdRCur6JrqDlAh17kpT
9e6ignmlNWJHlGz4yOQBwe1Ugvhpj/GMF1979+sZoCEK3ITXP0cvVaAIPbnIt1QO
51xOagEoY8vFIVwwQrp2REORO2ktaXp0yjsnAzgFK4/0Yb5hf1zoZzGjzdOQn7A5
WBYQlfvA9240yN+2YQb8PZ5WHgGeZCt1gXljhuk1OSuiwH7YpYKl9LRxyZPW2MeQ
0RK0R6+o1g2gWnzllWs4fdHRJ6JzZvgT9U3G+pqNoOPUvNNNs0GKcrmRNB1SKtaf
ux5iWWFRYTqj1phkYkPql7JT9JP9CFQaI/D0q4XtPe5Dsk2izw7qaR7NSW0bjxs1
ZpCnJIPugor5Vaw87snWtNgGBPdFXZD4UPggA/MeEz7sXBLzefgVp6R2tnv7AD7E
ur6Y6PPPjHiPkShzakPzu0Azq23T0MnnxKGNo8RMLUjHo5YkGeDb3CGH+/V1u+xx
WWElPRMGeIWa7oOaguOlyDo3x44gG/D1ZyiUMGnHQMWXI/GJNAEVBouCwA8UTddU
KWFmsDrE9UxFgAwJNluM022TXDjmb+lyhp+pxJJDZTCC+bHJd+hUgPvbxMVp7wYU
JUSWLRIiChHcz8KMmR+u1vJP+7y9nd2WrvwsM59+7CPLQi2R+fH/QNcpwYLSTJ4l
54WmISNfFy1qkVjf5DqFkJVb+jSBE/MLj56pfLJYQeyZQAsLc/imIjVyeM08RYn7
GyVWjDdex6XJdGgkJDmM978jEhYC41yYtWYVfUxC1AF1orURurWF/mXnhBOufBC0
Ym805zYq5tV6fqMg2w0mOvtdwgaE9Ap+ced5dOLQVjtU2CJ3H5iALUBIqa1UMqWY
YH5c3rlfKTANGrYhPK8vo0gXrWLEv1V2pbLSt5AwcwYS9dhaAuyjtrqqgKyfW46N
ApA91EkGy9fwZqaEiV2qjTe8I+EONQhv6/uy37DOo117TUMvg81a8M93gkwis0Tv
9hYRSXmDZlLOC6EmeXfsBx3FXrUiqHLoUHprroDaJMdAKCHQTQf0ic52tIt9XO+M
bDZtuoUuvlW4bD1tNy1+vqGSncPHc5QdsLZy3CDqjlgwVkk6KgOdyfSSLb+Kbwr6
Z6UEvizmL8iFaAiY94mdH8gojtYuZF8hMT/2qnQngkcON2HVkiRJDWxGXT3BanYi
Ixde0qumY5EkGT/nbiUeMRoGrbNTIFOwf4iy0RM0VkrVqbsGdSAAcORiIu04fXTY
JZ/QoajbxNbkc6iUjdAW/zNpgrMAjRpT87VXdBbxG+435FTO1XW8lvouI3n6HgZ3
xiPm1kNSsrTW0IuvvDgg9l2z5EoeG7q81V5pZiexpS0XMURgUTN0Xvbf08O+fe8B
bde75D5WuNt9+af3k+EzD5Tk9QR7dtdWzxOVZU0DGVa6E+D58s/j8+9oxDqXDoEk
6UTP4Ic5HnguJ22FgqwcTuLhl7xYivMpDbjHUiwOHy4YR6Ff58sRFWTxWQ5goEsO
xTYQG+KQSZQqkfLuaoEPrqjiH3YztgmQ50ocyCRulmn3Jz28PsINstkshp7lt1vE
WyK7GuTKydLL47wST0j+ws/Iu1Q0qXpjSiebVP+NCmQN9qn5gTmE6VXtm5Zd/oC6
rD9MwmVR6CZlQy25GbUi3IA8tNvDKKOIrKHwlBmIJ5g4YqS3DKV6Mcb0TItoNYb3
VCh+WxJHs15XoSg80gUVteuoelP8/sY9kvORFtVdZoPPlvXNZmHZo4t0gQLT9kRP
Wc+05EFg453MyhV02deQMoiYn5ajurLKqvyvSfy1A04TEN3lN6T30eoHosKILYhV
Rw1+znvlTX2hIyhtsYREmVKGGqEVEuJ5TucH3MvV5mFatXzdgpZ+28yncS/FSC+9
jitnHhh1Vmm6sK7rHdysTLCiVT+9reLmtjI98nmRwvJvs1o+LroRLs1qB/alo51p
RomaACmttC3hymepTkVrZUs42RIjZ61xMwLcR9G3Q44QZ/R80qGEIZAVqaCnzgWL
ni0EfCbZN67V5nvfZQg4sbo2+vfUDPEubplOGmvnqYJ67Pe+QaOFFhDeza8F7BIQ
GS+CQRWIemKSAaQJ8CXOeXPOecCgw9paAhdFJSid60Wcwuod0ZhgQA3qRUSF11ue
Q6r3i4ZxBM1zbF6q03jK6zkCslIwZD05wxOJZ8YlSuxSYD2wqrwTEKKKLrJITnX1
c2oNY6dS9X0AnXobPSWZrAIUOQnedn4oon1UqFTIAp8Bu6sZl7zgo2fUgO1Ds8ZH
PBRqKLYSGw5/PuhSoSsRB8NwQABAF5n1wsk+F9FAbT15SDaA/SNbOJHoV9pw0Kkd
Q5rnHSCFZ9z+Ay2pi8HyCyBBcN4I1vUhXtgXXdM0zRzUIKlvy+0VDZ6NyRBSqo1I
U0R5Fml7u0to8NnN+VMU6ShOygbnMIB67tBQmWnuMZ5M6cvyTAY8cVdJeTyFaRiD
sOSUcRjbwrm+Sdl5bvoLcnmze1L6H+md74y3C1AW1RshtvfnY6a/gN22Q9FgH6wy
xhXJmIgOI6AE01nOqrHmdk64k75moilnIp1SwRU55FJzFH/PVcw9knba5C9V9OuZ
cw3hP0UcgCzv2hKeDjx04YgddsXONQZvjK+sg9XXeeeOEIJwuBUgzxzgRCl+xEL7
oK7kVAMC3/ZwB1alxIYGQQDWj44DrI+LbjfJEcE889N57H/eG/nojnQxBye32new
nBFnnZo0GoJqzMcX+QYfZ7xPzUcT9SaisOXZWlXcGWYWc7NDSZfwovim/PT/ephR
WBDehv1HEIeqxtl5z7bZjZtVrDA6ZczbjHyYdqyp/Z2bwPy/MDxJWFkjb+sUskkv
fBmXMXrlnKoXZmvwIi1XLFXpefj6sYTyPr3yKwOILMZEzf69MUknUO+F2Ye9woDd
iExEwGsi22isSL/JwzoUgm99VGObPm1b66oadBPWNo/nO1/cpIkxEd/W6Cji+Z5v
SDePCTHJ+m/P37mPxc20V2zSiJZQSUDQgM+/LJ3DTkd89xqqddlQ3BaJ+BCrpR3D
tsaGm7X0ODuSgCz5vzUjr9zq/J7Dl7sDSP0n0lmdigstnp5djlkYH8Wc4XWBHErB
58uED11khEQMma0/ao4hQ1BNgFOqdNxFtxOvQfifis7N21S9AdWWAt7sX+Tqky7V
vJ+XhHu9zCte5iTCBVABOlNXKE9R52jy+wYOXwaVF7EK+axIrTUBkjXnenF5S2zJ
DFnF8p6rTsEcWWgaarnG250ah98P2ZEFJxGv9cmp3NAVWK3jaX3gZuputV8blwNe
wi1E5E8bYbWWemUP3YBGv7zMHR8ru5XxeiAlbU16Ssk5cg32UFUmnf3WxWOOrawy
cRAuFWfmK+9OTxRq+AzuJN/z2o85ZPorAVgu1X1FOgMnPeCWfoihM+xSiTPZPCzj
/NyHmOkfmXPWKVO1DYBO40hpbQfaiHztrAD2vb4eJPFQX/FtXhYi6ZcN+ba9hqwG
F7tCX976tANnriIk2kJUw26b7Qx3xolXhaXLngj7jodBIIEDTRYoxd1N6GhrwW1u
lITSlGrrWYPqf8zZ8UzcRZs6CSxl54nY/MJeLHkOAGBfHwBSJxTQdK8zAxIevqYm
L/unT4NyncgvRpQPm7ye+xL7hXCVJG6HKVfI+29s6N/5qbQ+l6thtvw5yS3PfYNX
+Vy37xVaAHJSltBrK9bnSB+zb3pa22gNGIMPNS2NWJ4tajUhfjh7+aqiJwPS92Uw
5AJQd6zV/ejNhCvw1tzpJzOmltqBYEiwc5OkPAbujLB50Si2DKWE3VQPR3OqLPJ5
BPq9KROsSlodkl+8HzEHVLoYJvJSsoQrWvjDy0KENPS8XXZawEELR6irquvFg+MD
d81+2mggL/eqWDUiDs3aIuT8MYjfLT1Pur+x2RJ7LVQtWLBPy+QwK1clhIrLnAkc
JwTnYTOXrCoXS2weJ1PoapOGfidVxcrUwvgiW5AAOBdM8DSIMe8IJz1lm69+BWcS
/PjbZc4wiaxRiEVI2rul80HVKmRjgyhcNa2YxNytQ3aVN8or1cl04yrSp2jG5wcT
hYs0d3p7OACqY/irFyM62veJfzxsKO1xknyJFjWL7D7zq1tgTlN0MhQH1bPhT8Xm
QEKC1Fy/jhQKBJGNrKsWzLIyjiTQ7IAMJk74g1Yovkb9GsBG7Aj07F6fqKMFLDsm
oHzd45feLbo6UXcZFdl4e1PDTJF0aZrL41wuaN5PV2eJAWpCwsWg/6JWOtC/4pQC
IWQ61JvJAVTYKo5Ld/rjA7jTnptivET7nLMKKBOnTI9zCAjL7XKSBH4/puqYzxB5
QLrajmMneWGHxojEcyZH6G/9E2kfC2RybC1YfPeu58SEBVfJJkDNO+pxmUJL+Z1K
UsBL1Ol3HYpLQ7m9Me3FSLUdLTqXPAvFrS+wMfDfmPfR8QiHnyEAi+71b5rTwFWI
YO5gp+jqsypX/tRFf4IsffqHjTadIYF2/HedDzzjNFCrFPzZVwfawnsXBM8swVjg
Td24zdnwZisgUTXnnRBMxTXPB4sFqLkHGwc4b8ueuBveoWzLKF02VeI7bYjd6doq
E7803VvPG/LsFoMT8+u6UEEOAd2K5N9nh1+Ws0YZWRThAuswxrkVq0aTClhyZXET
S1y/wrvF+n87pCA27u+FvAhAlY8mP+ex3iqsmFE6rtZxZnf/Q5qRq9wv6cLPYYkb
H5CC11JFda0R/u8WJjRM6So5O32wutd60CvxPYTAvzIpofrimoUyu6WplPv50BoU
agKf4tzlETBJ4citGyxSdtm3Xyj+2UiEnZp3oXyQRH/m6JMd0u66yyYjOgpNK+Qg
YAgNtaIt3zhsSOToFd4vWZKeU8KgUM5LAJ3bHP/Y/NUJFz34jQZqK5/36U1xsnyd
t9c853lYXoQvGlw8dIqHr48TKw2/nBfQSWeH+UtnGLOgVPBoZtomiE4JoIydRz5K
XYwJXdXcUsix8YZNbGEVMjxAvLHMOo8fAJiucl7/2jpcpWeAb0d1nQdiAbNsqclN
Pn6h/3NUjLpRz/uwYlz2SFbAbZRPy/bh6Imz0RJzszozRjv5QpUqaQt6MwK0aK/E
0XXa/W1oxAZ4E4WM5tJ4Q6eS/RmS2aJUQ1O1ZdAGPgz2CytfafFiR+vpWbaFEgy4
CmGym46j1QjIY4/tOzbP4UPob+85ZYTOoaDv8Bdfp3+ATZnhahdtVpF8Jf9hQlS+
iSeg8ikMcMCbmsVhCQ+IwKXwE4MIP7kpmw+qUtNAUQNPSk1llFPSuu7/bnEwwSOR
U3X0buQ8yzz8JETZvRIJ0ioRODRjehM7lFIXWlkwd+XjX4XqNpXqCwbDl1/sKHoF
A44lCWKKJi0fAZIRH29I13DjA4BGlho2IRqMtmOGoK35VZXPCqnIvuZXm+U4hLg7
mtdl6+f/HOwi5OX6UCS7yDaVBS5xPKaTCGZzMcDF005JpBsdKgljtCBkW4vqjoo0
AOcVjoHKBvfyM6PMxbd3dMloWL2aySGObMGhyJvRVJ07H2bzTA85JACOFJbf4iOB
LdmGCN+87fKDZzazcdMuluIk10PcNAIAJF2LNM5ZVYqYDP+eUpigULCNR97yJ8L0
Psl3OD8UZ+tMafoQC1IhE8vWMLlzvP2MZxKNNOiMyj4VSycRVMVLmAAIEZuMHkwu
A7ysyOO3E7X5ImSHNq2HYUHYnxsnfY2wR0HVpWfE3eCdOYY/421+xsuG25jJFFrl
gxwUn5meqVI+Cjf+Ceg/Qb40xB+fxBU+8dcrzCJfgjkFv9tazg9cJdlUKQoadYxz
M0UfOmRC84awdKiuQvoQ7iORF0po+kbpWE7FWLVUnqhwSuQHpVTzZaw9SjnUXxTq
zQddNTLu310djdNGRwstP57g5E9RkIBAnCazFpagqy15yX8+ijvIWEvN4W8lsOxA
Sj9Qa3x8/cVdorc2TjllAB4GfqfJ8rdK2QWHBFHgzBNRDKOGHJnnubT5UyTwzMNS
SJrVr3PJHYFQtRnN1Qr+MvvP3GV8xbohJ/p6HUikWb5gQt7aDKG4bY6iYwiM8OjM
PQiVTmmqHTPv7VSL5fS+90Xi0BCwb6svZaEbKDCsPCor/s4oo4kv1S59PjEZLD56
fleAY1fWdzxRWxDgTAD1UlWxLBVPCbq8VjwzNxidBSJI5jYQyXfPVgLrvrbbVZBj
6OQI4nDJmzEw7zyyPO+oXgnmW6qWXbvibO+8r6a+dpxCIudfrAupBVxiYfwSV1SR
B/GszMikXPyDnDK7/kCAndacroqcTXZmzhLw8Sv2HMI4ME7u4qHUus4LJTt8Wj+K
DAMnzt6gO36rLMrt/Vq7Yl4ThcYnPhXjix/gY9Cep32ZtO94pTAw93dKUE3pSJMG
TI8nyepEkKZDIiff8StZD95L0nEltOAJyPkoRXXudz/T6eHF2WNRj3OEMZhxeTqA
lQVzTh643vvnY07rtJAywTpDW4/rZ6zfBwR4tpAq+9vxEj/qbosaG5u8AcyhesHe
lgW2ru2Jg8tuuEEhYO2JsVTEi5cyIz4Gw4bsr5KB3lQYKVRir0lPcEAjAxSlmdIQ
PerUSNqKCP3eoJVgKwMXyDYrl+0HfngejwKgEbPwDxVnQanpkJ+fuPEub7DBhF1K
76DZ9B0sn4mI5rmFvYZCr9JUDbXkY0NRf9VU+BQQpoX/dw6gn6sA2p3G1ZVXKO29
LfSqef1M9fvlHvRomsxD+nUtZnBSfpZWaV7y4DO7JVDpRLFtakgoQP2vIIq1DjbJ
1CmHVdzc8Lo0qa1ghzoujtA7MdhnUZ2HkTUeViovakB43jV5l/SScoZrlhub4WCC
MrPKLRGNBjW7ziFKls1lzd853Hnkd/afdKpI1JQthTh0VId9ei3esfV3G2/TAk99
4cqS3o2TWV+M13J70FDuSUnZBUZTQhqnnAs3Tehw4qXlwALU3wXkRDWPtbhZVkuG
HlOxEtFyBtq5wUwY24eldw+BfL1yVF0e0bb7uvQORAAtsR3oBKEAaykiKFnD2NTL
Sg2iCSGOAA0IoT4cxcIxEk4oZ1raXIyHyNTeFWxoj0M96/5yTNj2OiQR2ku7hvg7
vgEosZzuTnS1CRL/u3erOuTdKHfNYWJjNHAOE4nb8jhAQ4rErS+Yt+ymUTbw2YL2
OhNBT5ZFQ4Qo09xZofnFo/5ymUjxQYRHECoCZGBsadq92Y+5BvOS+Y5Ty58GbAox
Y05dbHmRvolfWs+/Qi2JzGZ8VainZQS2/o9L95WEr9A5DLjfzw79zT2bRV5zvsAb
wNujUGyjjy3d5kPs+22uLTTNdV0HryL7pd9NbiuQLTiZCUmNtSA0e8vZnXY9KKUx
QLymX26va28MviRAuzgsNMHlwFUepYXgWNjiZOM/yO8qpLwgsqOn/RtO23hpxVJX
iMe2nNMAXy4gK+2Nftvrr8TqQb0BpVejuQISngJcv4pXnsI43iFhIm4WQ1TYilho
G5g8CCJC3eT+fSNHh3TGzZQvEzOhI1fY16cdn0h4ITmbp0s8Fr4hDPhHOdswoGrc
1+emkneqCHV9m2TSss4yF3m7+7ik0IDEp3kZ3RWDsa7843oLLIGttjNfLVmf+EWt
69JQd+YgIN4nOlxJnwkG26PFLAX3Bc9O1bDTo+KPZvGJCsht0sRbaa6lL071UB2q
zd7aPDRK8Q4lOppwe4NZRIkKeG6Jge3UJMVYLRt3zGbaRHHq2bSAH1kgKV32CfXC
X0lbD+ln4nZZrMnp5XE4XFjZNtW27ZQr3RIDzX6ZnXHMDc3ju/CsFYS0dP9RuMca
oVds6LZfMQi5ZHY24UyOTN24484PWNEODEs59bIqaOzjLRaQgHpU7Lm65MxvZO4p
k48f0jZiO4CAjnOfdWVHtYQKXQJ0CjcDJsslS1dUPQoUcinkuYJeoqxqS97Px1rf
ENj+kgXT2p3Q/T31AOTHA0gu9D/MUDKI+UXNJ8RlNncZAhUKo53Lmz8eaEcDAFsq
m9HyRTh6swNjakK4HN8JpWwxGgJhkik/jKeOQJusM7iT5VclRnjINqwSc9cHdHXS
dLs3S7gZDBrMupLlPyriDmUzcH62CckFQkUy2rdLRqVw4pGQ7Z7clBCoURYbAmJk
RMc/W3escZ9gszxyqNDMsTDyEOR9l4PLodfQV9+Q/wkIi6dcfVYg1dTJvk7NIcQI
g9P8a0jQ3EIZrFWqgN6ylcfpOVLKJsy+qi7MRYueCsXiUB6nLbMK6+oMPpDdxT96
zhwNBJE9ws1cuAenMIR+rKsxeplN2OIC8J7Vmiyn8Kmb75f37GM5JqZ5Q+EpI8/B
An2jcWUz67j99/7UBE0NGmukRoXUmEJdjDYbXOEdPwBSMSXcZxTCPzhYfM7Y3/Fq
5pfAIsHfieU7On9vct3fRYu0yPUcEEF0FMvbaJgExAkeowotlXeFeIyS1xA8PCCC
Su3BfrHoNWd31SgZQWRQ6tyOfMT+Bi5TRgMhhe9BQBQVZVs8/7UCO/wLlNNLE6Yr
mZoO7IUxRS9qbXk37vAOCsTdbgc4sTeRC/PzTErqb+ESM7N92YAYVP1ba94U17+x
+8eRJ/N527OHX70gi8CcJvSnay/ppN2p0r97iCJAnA8uGoE1nvCXYbF4s5VGBgZp
mbleb8fOijzCkJNpenGuAFuhSImCIuZn/d5NjLMTJePwM5cnT8lGgd6AEmrnEx/u
hbCRTRAwP8sIY9XZLVJ4FGHoxaRmtUTHedhJXWrCOWocZdMTkl2zekPH4PHjD3Ib
XPRXcCDvYa4eIEJStlFouU+EPOoyoZJj45BD5sywPq1vLe/yDT8VkMesO7RKHfiA
Tb1zq7lQhbM/5gnqtaEU+kDaZF4xi5l2anpma5CjYSPaqJp2hU5LYGKdpxKMKp/o
9sBJUSwprPjh7OaabjmPSXUZyZuYZBp+N1AGHyb5S29B90WpJDHcHdwJHHPpJqKV
kbPyiO/ERAwy0jkQ4cpy9q8K0UNff8IY/h5hdCcp4EDIGlqNfsdk2ypfqfSSDhT3
i2NUBLO8SPPYM7bKy6O3yCxvtMYyLagtYSiIzsPGmyf0XyIaWT0mn8m/S/Jo1/Mt
OtIa+o/I8spz2i6fi6eK4KIYJ+FVu+M8sErsVO805Z3R2UchLEUThs2jbqP7sY7h
ebdO59g4Sg/Lld54JHkQP7FxJJRtdYn5hqaDc8Hd4w1qPu0DaITJuRe4WhogJodr
jfo5eBulsJvlQzf80g6sqt4CzupnzyxLF6yehsvEX5ylZHkriVkzk60Dd4pa3rLQ
/fP9nnHI7PrWC6P1Og0ns7j+oZFiAEyylDmaCckpzl5tQrSvGPqRsgucOAwPEKRX
FCTJ1IZK2RFcsOhsW2zM7gAsdCD/Z7uBYPKQL/nLfJyaA68sVljZOJN+Tjqzkrxu
Zf0r0xEOBkQOJHSZ88r2iTZmBeL1WtYkf7bpW+0FwvjnUt243xZt9jeKrUyneXOp
p1PitDS5zdNyWdpvD4nNiCWScPFisHs65UB8XCZbX+i5knQj2XCZ/ekIkzT51oiE
5lxS6U8xRbaqkR8qyGBJPzm82DprsrRyWU69rBBZj4GVHFCKyChZnxbP6fTjvdtF
uGFfA/jX2NgmCoEkQf2yWmUy9iMqHs7AF9D2YaCZGU3fVF5ZgVjBfF/raBmlB875
rBYspwH4T9JjS32fo+J+cpIxErOtvJA5+eo9mPBNZiPEkKxw0MDVZIRUjZF+2dQg
sOfTCLTx3WkVk8wx9SLN0x8c7eSKS7WEjyxpX/vLNCUl0eTI2jAkveiwa7B/ivi2
gnXsbdGV83W2cv1y3MWExGvvmfSPhrmg0z9roONHZYBYdIFLPod89eYr8LEN5x/W
GH0hk1Vu6ftw43aQcg/Qx/lGWVXT1Yn+1ufaXZuNXhWjUDawWktio1gYlAoyioAZ
YyC8rmzw+BhTkFrJZYZ7Nr9cCGZ50rjsS0qwQ4LPW4rn6Ur3g9U6v3OmU5FJzJw4
Zy7aO2wwhfA4SRD2nRMgVBAHVwrZeFhaugD10k74ZGobnXCCLmjxljtm48oyboov
1bygQuec8SthN/mzpFKldHHyVFPqffodQi8BQwMhi+Dn34Gm6ZE4D1E1l7Khkkl9
Kzs66gx8MJil5wskNcI5HvdvQx0OLy4sfV51jyAHqDJzwyWpJHpbFJa2ro8USVhs
XHO06DEF5ySe4mMWNDiDTrzvTFU+/MwQf4kgl4AUkexJkkjDcdaQJ4xU8+Jx9opl
0wKqDXE24eyLozj7MJNaJ1fm+jXt9G4oOeBmE5PhAtLiDRm1B7EIkwY5M5/XAnmX
DoY+MhN6aQp+cqf6+oD6ieJG3q2ia3AtRBRyK/ey/Eo3bhsgq3jOPfAqtxmP6sQy
d7qtwdn0UN6GLIGVj+UFLt+1sFyeCBdoLpu41wO7/l+ndyvcaIpAipzspFeV8SXy
heVrN1/yDldM92ieYBEhXtnG2i4olyxaqWgSmnPvqlxowCNCoMTDPoOx4PFao0/Y
zEFQ1dJWrspFJtYeK6QKxhVKULPDmXrIj+QDhBKmKju6Vwe8sVzrdq5I/zhJnn/d
bbAYeWpAu6T81lzGXuZbMWrZJq2bXsDQWmNqnjtRUCPqpiDvEwaPqeO/9dKrg2Ok
wcx6Fj672Ew4mSF1MyDQA4LU4BjoeRCCKYQeEYx4r8zvtkfxsMjQMFAFB9PTISdf
7zXitsrRYsc14hFCTci7xrw/v6WXdQvFvk3hNYcLBJSo138bZ/Qd3nU+cfmVDikX
7Hjvm4yVgp5j4TEPovYzCeat8T0obktAIRLcSD4CmmYmOUQHlDDAM4wamGQV/Ik3
poa0/Y45GNdf+HO9lxBkaWXsKPHv0Oe+nimaPt+vx7N2B29NlQNomK9g4UxvTBEV
fdThDr82uhuzgqABzQw1/chWY5divDRzFCj9iGurLqIFDu+KlFMfYZco/B7+5h4g
q+e/0kaIm6E3tM5SFUueMg==
//pragma protect end_data_block
//pragma protect digest_block
p2LTFrT9gj0g76mRZ4bgIQAKx0I=
//pragma protect end_digest_block
//pragma protect end_protected
